conectix             0���pycs   Wi2k   @      @   (�?   ���t�F�nWw'�Kw�rΦ�                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������            
     ���m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%PDF-1.7
%����
1 0 obj
<</Type/Catalog/Pages 2 0 R/Lang(fr) /StructTreeRoot 21 0 R/MarkInfo<</Marked true>>/Metadata 144 0 R/ViewerPreferences 145 0 R>>
endobj
2 0 obj
<</Type/Pages/Count 3/Kids[ 3 0 R 14 0 R 18 0 R] >>
endobj
3 0 obj
<</Type/Page/Parent 2 0 R/Resources<</Font<</F1 5 0 R/F2 9 0 R>>/ExtGState<</GS7 7 0 R/GS8 8 0 R>>/ProcSet[/PDF/Text/ImageB/ImageC/ImageI] >>/MediaBox[ 0 0 612 792] /Contents 4 0 R/Group<</Type/Group/S/Transparency/CS/DeviceRGB>>/Tabs/S/StructParents 0>>
endobj
4 0 obj
<</Filter/FlateDecode/Length 2986>>
stream
x��Z[o�8~���G{1aEݵ�I;��t��؇�}`d��ַ��_��B�v�V��m�"��s��!ś��^���7�>��ͯz=�����8�L���;����'=��)_x"���������_�������՛�J�Hf�x,�����'S?�������!ss�9�Jݯ���~�߭g�`�Wf]�o��^�o�B�o���4^�?��Q�������/�W�@�߮�~DV?����e%�d�t!�����DOI/|�8U2J;i)�+S��q82�l$:�L���'4��D�H-�
��>��91+m�#���.p�����hoh��X�#A��E	���@-b�y��d5c�:�������v�J��ssP��n�u�
�@�qXb���ĉT݅��M�x�um��ژ�E�|E��k��N�xѬB�%����/4j�F,#z��|2�fZ�i_EN!9M]~)q޺4v@��(�a҇���|T�˅rr�hd,��W�`F�#*�F�-�`�] ���n7kKO�K�~D��#�3Z��C4Bo�i����J ������A�@�Ts���-����5��qH�#}8]@!A*U7N���?`(�^ς�y��S�&k�%��qȀ��nQd��8h�� R�4Ŀ~�K�I�y7�QA�A/ G���AmއKQߛ��!���Xy2�t��`H��GSJ��Sȩ?�G��a�p	�x�U�ښ�k����Hzt���k��2�*�I�eQ���)�=CXGskSdW�ƨq�i�' ;�^^�|Z�(��9��!��c��޷���ǘ�W��4��?�H"c=��]L���䂚���Ҍ���L�0I#��q"J�׼E׍-��S��z����E���������y�Z��5��v�����L�Q��6���lA�*�Su��ʉb$@���4Cƿ �i����7�z-�� �w$o�h8�Yr����\���@���5�[��B�v�ZJ%�5�8�*�y���2�^,$`V.�"�n��׳��R����J�����V#Sʿ?�t]?��({Ĺ �*�^����E쒋�\��#Į�� .�}��n�eHf_'�X-1DL�39�-��9S�9�b@�pAY��*��V��)�
��6�c���ҽx�"¯�R?�|��x�S!3�\���9��σ�$@�{�8�5�"�!dX?�H�qXDi��
���hHN���T�.x�p8�t�r�#��<��O�3��.DA�0}ͫ^�ﴽ�w����<�#���W�e͆_"qpDA9Z���XC�����QA=�j�̢��P ���ܩ�ۊnH�R�}] ����ɚݻ�h�/�t���oE9����5��Z5�@�vjlM�����y0U���j��YWm�[Z�C�a䪛1�6��0m0�).���I��d}@]@#*�Y�dl?w�8P���G}e���(�_OT�Y*��~1�:5��� �`ni����݆��Nu���Ҭ�hԒ�j��.J�f6d�G��zเ�PF݅f������t�Dr�P�6ۡ����`�5���ƂAykؕtw��خs��@�S�3��6�I�ϐdЈ�@��5�^�f��3#����5��Ջ�҄+U�1q<��um����O4����Q��M8v-��j���O������Vm��Y�A�7�bx���C�P�J� <���WA�˴]_��B�>���l�	�>�gl_õ��g8n����e��I{~Ʌ(U�2얁-�:�-���1��vL�]VS���F����=T4�71�Q�AG 8&k����Dն-*�R\��-�W���z��_0����;�J�&j^Ps�> ��̺܌I���H�TDA9����2u�7$�<7*A�o0m����=雊T��ޚ������Ӗ�N#	ow���še͖ǽ�h���]����D�HM0��WSh]9�A��wS%C���5�g����!K���Z��� �KE��.W�m��L[9����: ꜰ�@BB��z�$�>�Q����[Y�`�y�F9�]40�8N�n\BW��4u��m��NR��(��߇�ԙz2���(Aa�m��9�����BӮLW��[w���7G�^�z��cGѷ������G�Qp����`¤�H�i�
T6
�|p͋(j:/����<�^��Q �n�F#i�w\���!Aۖ}�t���j\|��!���?'��л��p<)H}�D}os�مx��2�j|J�8-u0�� �ͧ�ua�G$�j��Wn��a���E�F6��Yұ-�x�˜�>�4R�	�9CN�:���ҏ��#]��v�gA�v���D��a+Ŵ��z	�w�/��m�٭���� >�;O�w�ӇO�S�V<��On"�����5��|.�&J��ѳ�<OLS��GD���WQSE{�a��=�M')���ΙM�ۍ�1�>I�[d^+e3r#)ҌVϦG�2e9�M��U����G9y��xC�������I<Qx�.�����AxD!�I&�Wŗ�k�N�'H(�M��u_�)�f�)b�y��H�n|$=�E"�`�ѡӫʲ�N@教Q� }i�]�Cٷ�9�.��j/I"�����-2Ǻ���%2���A.���ME�2��1ϥ�3{�U��N2��&�qd���ΈYh>��t��(>0~��Tj��I<��LP��<MŠ�������ES+2o�		.� � ���46��>�����c��ڟ[`w�P��-;2g(�wEѰ2&dݍ=T��61�ۓ��4u���v��K{V��"�?Le�=��@���>hS[b�n�1rlzrPDh��0���!�V��b�~*�I�봻�Kz�r�(eI��w7E�qeK�C�*�*kT�J�K�+��yix�a�����^윸����X���s�#ҥN8f>(�e���u�
endstream
endobj
5 0 obj
<</Type/Font/Subtype/TrueType/Name/F1/BaseFont/BCDEEE+Calibri/Encoding/WinAnsiEncoding/FontDescriptor 6 0 R/FirstChar 32/LastChar 122/Widths 141 0 R>>
endobj
6 0 obj
<</Type/FontDescriptor/FontName/BCDEEE+Calibri/Flags 32/ItalicAngle 0/Ascent 750/Descent -250/CapHeight 750/AvgWidth 521/MaxWidth 1743/FontWeight 400/XHeight 250/StemV 52/FontBBox[ -503 -250 1240 750] /FontFile2 139 0 R>>
endobj
7 0 obj
<</Type/ExtGState/BM/Normal/ca 1>>
endobj
8 0 obj
<</Type/ExtGState/BM/Normal/CA 1>>
endobj
9 0 obj
<</Type/Font/Subtype/Type0/BaseFont/BCDFEE+Calibri/Encoding/Identity-H/DescendantFonts 10 0 R/ToUnicode 138 0 R>>
endobj
10 0 obj
[ 11 0 R] 
endobj
11 0 obj
<</BaseFont/BCDFEE+Calibri/Subtype/CIDFontType2/Type/Font/CIDToGIDMap/Identity/DW 1000/CIDSystemInfo 12 0 R/FontDescriptor 13 0 R/W 140 0 R>>
endobj
12 0 obj
<</Ordering(Identity) /Registry(Adobe) /Supplement 0>>
endobj
13 0 obj
<</Type/FontDescriptor/FontName/BCDFEE+Calibri/Flags 32/ItalicAngle 0/Ascent 750/Descent -250/CapHeight 750/AvgWidth 521/MaxWidth 1743/FontWeight 400/XHeight 250/StemV 52/FontBBox[ -503 -250 1240 750] /FontFile2 139 0 R>>
endobj
14 0 obj
<</Type/Page/Parent 2 0 R/Resources<</Font<</F1 5 0 R/F3 16 0 R>>/ExtGState<</GS7 7 0 R/GS8 8 0 R>>/ProcSet[/PDF/Text/ImageB/ImageC/ImageI] >>/MediaBox[ 0 0 612 792] /Contents 15 0 R/Group<</Type/Group/S/Transparency/CS/DeviceRGB>>/Tabs/S/StructParents 1>>
endobj
15 0 obj
<</Filter/FlateDecode/Length 2751>>
stream
x���]o�6���?��^4������t�N������,�Z;�W�����=�P�儔�l '�M����yϡ�������w_����w���-��_�?��~�������|�ɸ`>��w�	V��W_��v�W?�]_��'g<��-��8��g��"�?�N���ݧۄ�$쓭�Y�>�t}�����<���M8��r�S�o�L�|��r����v�[��o��Ӿް�����g�r������#��_�Wo�7yI4�7h���yG�����O,��r��F��4�qʽ(}1"{E��?fܻ<8����e�'L�{5]o���0��> ?��4%�'��,�2�v�>�؊�tƪ+�I����|��9nl��
�x�F.2����l�
�(���a����]�
;���`���h�Ws�#�Z�H��ó� �鬩�R2�Mo-�x� �0j��4���lr�� �`��+u�sB��#�j�D��r7�H˛ d�p�LgO%bY���Mb�U=��YVϹ?#DMjɰ]�Һ@�sP͢��c�$�;�݈��X:"�O�M�����<��pЩ+�u�s���O�%`���p+G��� �-%�ǀ�4�BȖ؂����9�O0�Uސ6+�lq*�
�\a�yȥ��^�ڌA(��;x�kso@&s�s�q/�9��3��Y788����d�
�"`3V|����f�Y] �&@|A�dO�%���̌q�m� ��3[�h:��LS_�^�)l�rM��9�S���uްJ"[��~�~B��r~�ܯ����M+���&-��LWF�ɰ���vg�~�f�=έ͡�ػ�UQ��f2LW�J78'\j�1��.�$�ܖ(�m @))���b=�ьa����;@u�J��iM[k����D�皙�t
��<�vtNp�w���'�8E
'�n[��)4�wk_ �$�OH$��LQo��۪!R��'~JE�}� mj)�cQdm"M �2T�ϽxLL�)x�rT��9�S�ы����M�Q��zCjJ��ۡ�Vk�Z"r�$�*'�zO�J�k���Tjm�=�)��K#k3i"��A
�l\>�?%wo�"q_x�ax. 5tt~�b��N�W���*�GUI�E)�S�n󺤴U!55j�OI�Jnl^�c����5A��9�Q<��|R�ɺu���	����k�rx�o��!a�T]�	�ƛ������, p���|�Gݶ)ܦ+$�.�����` M��[�a��U�����R�֭U�nxN��w�a,wM�|�X����h�S��+V!r�g��(	�[*�e����V��*� '�&�t�]���_T��Z��n�:6u�s¦�#%�����Z����v�NIS̀�u1mJ�b0��*�>�}�k��c~떕�㜷o)S�Ӯ�r�T�$���ڴ�ppe��4���S
Uº�ji�����F�TX��|�a��T���3Th���8բ����RAY��cYS��lͣ���rUAJ4���S��Ui��O}G���ן���-ۢ�!����i���+�@T�,���b߮lA�մ��G�T�|�M�Jj�����5A��Ua�k�F��R�
\�*��0��H��$��
42��	CU� �bӪ����jaD������;Z��B�	aȇ���=`F��<����SBZ]��c�`눘Hr����d4ҝR�
\�0�𜀮��t3�t�@b��B�p�V/�u�� 8 _��)� 	���R�U��+`�6�⽔[�;�1we�D�]��)U���������ƫ��7R��ZEH���f������$*Zm5F�D�&�c΃�X
}����a},��!4,��H�ִ�pqe�D_�)E���9��	���H`%�P�" ����Jl�R	j��[���a2�N����o�\�
-�^��ƪC��&��hF�ŰaS��Sb�&��+'���R]�8��p����Z�i��A U�J�
����ƒ��
ZSv�iK�`���J� .F5�d�
���I���A��T�}�m�{<�6�&f\�<\�}Ŕ�Y���i��i}G]b�>ߵц���j�C�}��:c�bz�l�+7G�m�V���ښd�|��/�b��^�|�vxN��wt$�	>L��A$�A.6e�RQ��T7��Vm�-����aK�^2�]WXr��L9YB�ki�Ml��w<��t��BW�N;<�:����'��V5�kh%�"o�{Lm�������#�o(���U��
Nb��n��f�YaP[nm�Mh��rB��:��Rg]Y9��p��ǘ.�V�R�z�]U�%5nW0�s�nY ݟV�/�j��3|���79��g�����6�����7�����_�)�ȕ���	���Fl�RE�.�5e
��m-����d˚�eխ�}ʷ[v~kòZ�'�*)nJ�Q�ѯ��6!�ʹq����\�ʸ�F�_m?�zr�.!�ͺ�pXW3ko��h�>���H�tD٨���Пa6aP�����9�W?#�t��s�I�vY����>���!-Fa��ZK��D�+w�a|4��S�r�+w���iCd�e_,��R�Z,�^��vudN;���/��Ee��&�L�������R�&��=H���7q���%.��XO��E���vx.�6t4�!ה����5
S�2Nk�k8�Q:���,Z�*�	q��rPO��&gI�j��*&D~ӯ���{y��a�p�?��
endstream
endobj
16 0 obj
<</Type/Font/Subtype/TrueType/Name/F3/BaseFont/BCDGEE+ArialMT/Encoding/WinAnsiEncoding/FontDescriptor 17 0 R/FirstChar 32/LastChar 32/Widths 142 0 R>>
endobj
17 0 obj
<</Type/FontDescriptor/FontName/BCDGEE+ArialMT/Flags 32/ItalicAngle 0/Ascent 905/Descent -210/CapHeight 728/AvgWidth 441/MaxWidth 2665/FontWeight 400/XHeight 250/Leading 33/StemV 44/FontBBox[ -665 -210 2000 728] /FontFile2 143 0 R>>
endobj
18 0 obj
<</Type/Page/Parent 2 0 R/Resources<</Font<</F1 5 0 R/F3 16 0 R>>/ExtGState<</GS7 7 0 R/GS8 8 0 R>>/ProcSet[/PDF/Text/ImageB/ImageC/ImageI] >>/MediaBox[ 0 0 612 792] /Contents 19 0 R/Group<</Type/Group/S/Transparency/CS/DeviceRGB>>/Tabs/S/StructParents 2>>
endobj
19 0 obj
<</Filter/FlateDecode/Length 478>>
stream
x���Qk�0����(�H�k9P��$+�È��4Wv��Y��ߝ�e4ݠ���������w0Y����r�ab�I�X�'�%������ǑH]S����j�Ao���;pqt[���)SQ@�ƑD� 	U�VYJ�T�P?��n����U��.� ����y`�4�_��G�����_���~��Ru�7���:zKc�(�3�
-�wm�s<g0�$gk��݆K�vz��=�WlX[�4�K�6�lyR��%����`��>��0T��2c�3}��%�0�u�QG%zÓ���G���k�چK�L:^c��J���'��%������X��?��/����.���Bs����x��7.�i�{���R�D�!���{��`�	����xz��C��=�!��6�(8�<�<��`�dG3 �m���׃��8N	N��a�e��]�W:6�Ł(����+�罼"��a;8�B.X�
endstream
endobj
20 0 obj
<</Author(BiServ) /Creator(�� M i c r o s o f t �   W o r d   2 0 1 6) /CreationDate(D:20260107084912+01'00') /ModDate(D:20260107084912+01'00') /Producer(�� M i c r o s o f t �   W o r d   2 0 1 6) >>
endobj
28 0 obj
<</Type/ObjStm/N 115/First 936/Filter/FlateDecode/Length 1725>>
stream
x��YMo�8���q�$���~�E� H
���M����*h����ZRIqM`/�h���f4�0�e�3͙lo��q-�L��IɄ�L�5L�J[&S�c�2�=��-�����WLqfn3�rǔe��7͜��3�%�-��A9,�b(�i0�d�A�8�kƅ����2���I#Nan �
��؉!�^1`�Kl��A��������8'�A�,-P�Ay�B?>v�زEF$�d>�(�
;��S�c���e5>=g�J���r����bq���X�S����t�R�1RO��-�;�ԡ6
c�Axϰ��؜G���P �H�2x���55�R(�&�
���'��#��n�bFO��f�� +��~yK��<A�r�1��>%�=�j\ Y�E8�P��ʋ�kL���3s�l,U��$D=�pl�cfG�&6yDp"�G:9v�[p��6�_��D��*-.�P��@�����Q��������6����撘E\#�8�㨭v�X�U��KMK�×fXS�Zb>QLA�� ���b<*�XL �Z���\�A�<{֜�,-�h.������]sy�?^^�u���Ϭ��&��ϟ>�!��qz�<=D��O1����C��!���5寨?� @�!Oc�����
9�Q��?W���cܻ$��/Ȩ���Õ��\U�p�,���}��Յ�\S�>��y�j�-D��*�:�5y�v�/D���T
x]��xM[�ZZlǰ,�*���f�,��r;�eW�ͨ X�����aY�U�36 vy�� 8-�cXp���@5z���� 8-�cX�0�Dge ��'Ң�e���g�g'Ң�E�U����\��\��DZt��r�Jt.؜�ۜ+؜H���\%:�����N�E�N'�D�ӹ�����ɴ�|��d��|p:�w:_p:��/:���N��N�N'Ӣ�E��U����|��|��dZt��t�Jt�h!��g�A��:��&q��F��@���Z?��UZ{��,�*�Qw*��{5��A��7�˂� ���<�{�.[���$.�J�������y��TZ���,�:!rA���Z��3B�E�uB�.��{ 5?WA�E�u�E�Aj��A�Pg�(�N��(T��Bj���Q�P�	Q�:���^=��²G�d`	��~(��X�-������A�Ԑ:�WK�C�V0�O�a&[8A'���E�{�c���tό�$�7�����n|o�oc�g|m�x4��/�G��T��F:��f���}��-%6��?�ݟl��d6ݠ�S�_D�����z��v���o�C�J$��ea{,� ���}��<�Wt���0�
���5}'�`��ﺋ�?4�]�q�gs��5���co8����Y�����d�������9�?�w���'�����\vW��m�����b��w�����B���3l�~�����.������׾�v�3}�p�uyh>n���d��'�W��]3���n{�����f��o�lo����p�5oy󲿧U_�n�}���a��)9{�����L���P��nӺ�m�a�����G�L�!1������n��<o�λ����6on�;G�̼�1o(�O�����9?�-OH����~�ʼ|]��-ߡ��'K���T�N�Zz��9��ɿ|}O�
endstream
endobj
44 0 obj
<</O/List/ListNumbering/Decimal>>
endobj
138 0 obj
<</Filter/FlateDecode/Length 356>>
stream
x�}�Mn�0�����t���ABH	)���i@̐"c���53$m��%�>�{�x~^Jݎ���:�ȚV���b��[��-�[5.�o�U���8#t�nz/M����h'����	<���`[}f�����x1�:�#�,c54�<W0m�v�v����x�0��i��0�J����4p'ci�N恮��\�F}V��d�x �"��Eů�k����bQS=�k���d[l��B$EH�r�$Z|1с(A�r�=QA��?�ql���g��~l�4,�E� I�N1��)��冈Ɩ��>$�usI�KlB���h�H8��%�?8�u��%ӈ����j���fv��7�U�m
endstream
endobj
139 0 obj
<</Filter/FlateDecode/Length 62811/Length1 157120>>
stream
x��}	XTG���{��Y�U��nl�w�i��J�7�E4����,jBb��jV�g�I�V#f����g�M2�d��&f2&���=]Jg�{�|�?}��[��έ�[U�ZQH�U������ �^�{Z^��Gf��kQ�瓦f���a��y�UQ��rqjh�WDg\Nd^S�b�s�⷇���k�]��}8��5sn��ڰ7�> ��SI���TV�8a��"oXֻ����H��[�|U�s����hގ�EU�tY҃��Q|ڂ�U��[3�!��j�W^s������;wa傚�M��X�xѲ�vڄ�xe��Kk���ޕh�(��K�c2����7;z�!�j!i|��y�o�����#�a,�'��Fl�BGI<��Ç��0"���;��އn"�"5m�E��b��ruS����d1o5F�Tf�eڤ���h��i&]3}J�[�Q��F`�:��&���m�A�p�h�y�s��)ś���F���}���0S>Uv�?@;ڧ��;����i�9�����c�5����4���놼����<�|U�+�0u�8�9Te�7w��N��E�+�8�BS�����=f߿h&ݤ?G:ͫ��n��c��1�n2�M�'�[u��8�뱐��6:���}�yݐ�����LwQ�ɴ]���15S�~�q�DE��)�nn<������4���4L?���ϣ��7h��ޫ�}Ch�>��;�]D�!���Q����~��'sm	��\C�7(ݴ�ڀE�'S?d�ɕS�d��0�#��{�<��c��^��?NCO�u\_��J�7i�o�e��T:O���	��o�gkguC�ik���Ж�Ο�/�Ē�Ҟ�WO��������1?�4SCG_��Fs��c~����e����*�L����[N|��J��H�O����_���|�/T�M4x��Bc�~�]E}�/�^TQ�X��6��b՛���g
�z�#~ �\�	�dm#9������zi�ȡ�ܓ���a^�x��nEЂ���i׊p�����Z4�մF2>c�1�=��LW�rʯ��4mm֜�wӹ���*w2�����/��r��=G.� �JLꮿFt?W3�yxp��8���
�b ��j[��~�ЗQ���2�:����B���0G��i
���-@0	�*�Y@�,sB�z�t�t�>��Ɖq��Q�v7��ޣt�v�3>��ڥ4H��;~R��O�j�S�8D�)4J+�~�x��
Q��h��];�& �I��;K���o���ڟ}tf�!��=���b�H���.��N��颶�H� ��f�ko�\��N��{���m'~FZЂ��-hAZЂ����m�3�2�9�п�9�(��/*?o�5�3��1���-hAZЂ��-hAZ�~?��S�AZЂ��-hAZЂ��-hA��c�b���@�
��v ^����4�L
�?P�c�ԝ�n��?�wЂ��-hAZЂ��-hAZЂ��-hAZЂ��-h�l����-Z�~g��ƿIJ����$��.8��Mf���Rw�M}�?��CETJ���F;i��O�20eh�ȔQ)�\g���s�s��|�E���dj5~O�8��e�%�NC�JD�E�28%QF�EY�\�܂(�(���7M��G�>f�M�z����4�u����I�'�>�D�����2�ߙ�� �.�����S�����o��t}�~�~@?�������]�^?��N���͠��i�OT�~��.��Zh"Z�D�H��dQ.f�y�^,b�X/���%��[��œ�)�I7��G&�)�j���L�S��j����+�E1�����p��CZ�1�~ݸ�ѻv�d�~���t�oUz�1g:���qcax�wҌc�~�����w�<�7�ɧy�AEmp�vj��W*��7m\�l�ŋ.�?c�����5�sfϚ9czy��S:uJ��I'�V<�h�����1�ѧ�:e���Æf��׷WFzWwGR|�-�f	1�tMP�Wa�ӗQ�3e�ƍ�'ӮJ8*�9*|N�
;��9+�bΎ%�(Y{\I7�t��6�(կ��������r���/��|W��w��m�0V$��P�Y�T���
g��pE]SAE>�5G���j�������(_/��f�k�0�֫`d�F���OO/���M.��������|!y�P#�s�l3]�l��ͩȌ�vUW����JTj���6�b2}�]���k>MB�k|}]��L�Oi����m.g�!B�]t�T<!�C$��b�0!_iB��B�/-M��7�A��X�崓������,�i2g��I�ȜF��V�&UAE�{E]��q��__���o�;}zFŜ�:ɕ5M��|�R�ϝ����y@�WV���0�x}Y�žxW.��)����^�J��/>�GU�Z���|�.gASE>7P�r�x���֏��8�;�*���%��d4y�k}�
{5�g��kO��0|e.oM�|J.���G�]�qG��v\iUX�<4���jv�L>-8����rG!Æ�e$����
;�b�K��T� ��獓Y���7ΞV���+M��dN�Y�Ų���&��/6�K��v��k`���@�:o�&�"pc԰��9Ne��X��ic��SLr�h���q��0�ܓ��or���[<�U\R�5�v`��vHq~6�|��l���03���F�-9��"���jj�n&=]Ne{�0�9�2ߤ�2�oN�+M��_�fE��V�a�b�sV��6gaSeKk㜦f��iqAE�H��&WQu�k�w��h��z�y�X*ť��Qn�K�W���M-��9�+��5��U�5�@�w�/ ëI�tʄS&d�)HX����x�5�&�a��Z>��	�j��g�e7r�W�b��*m��¾F.�+Pڂ�̹��"!#���� ���n�;��Y5�t��e��VaoF�)��E46���{�HS%QR��|h�,�.���끧ܻ3�߸�D�4�¤:�!�O
��r��+�k�(��%b��[��k4�4�h�8$����E�r�?G�s�"����"Q�a�M���+�Kv�kM�!�-���޴��Ұ�f �^_X&^n���(7V�ƪJ��xe�����2�KE�|a����F��P�
s��eH��u4���2�M��ʌ�j��8�H_H�4g�e�5ź��zx�fIahM��ǎ$nVƃ��W��UU��92k�_�v��`�7e��2IvKO������# ����/�szhY7�Hm��m��(��P*`t�U$ۂ��h�,�_�)i�)�U�:e��H���YӋ*�v���Ue��#1go��y$�[BK���i�{�|���G����Y�t��7=�__��^��nj�X;���e�����ҫ�[,'�1ߜ�U�߬M�4X�4ޅ7��.������.������^���D�B�5mo���R"�����1Yז,��a0�?�!���b�̷��13U�D�MN�k�K^��c%*�ږ�?f�\4�UN�Lv,�h*l�GԪ�����[��!$օ��A �_�dgE��GSQ�MK�c5���8��*�`2�gr�qT�l�S�pR)��B�b���q���;��l�)�l����j���>ˮH�g�*k��V��k���h�1:2�����\�1�8l}s䥪I�gVdb$b�b��#�����ÔQ5��*�Fr��Ҏ�H�����˂�dkd6�M?�1�era�-���MVE��$ŒL��%���bJ�W�S��.��1�첶ӧ�z�Ǩ_$����j����j{ۨ��;���x9�c�jOkOR69���>ek�G{��� �	~�:�5��W���?~�<d�ޣ!@)���j�V�u�Lg ����=J�@5��0���Ȼ9�sw�%��x��(q�g)ѨęJlPb��X��%V+�J��J�P�A��J,Sb���X��B%(Q��J�Wb�uJ�U�V�%���Rb��JT(1[�YJ�Tb�ӕ(W�L	��+1M	��JLUb�%JLVb�����iJ+1^�"%�)1V�B%
��W"O�\%�(�V"G��J���(%NQb�#��Vb�Ô��%+1H��JP"K��J�S���J�Q�����D��J�P¥Dw%Ҕp*�P"U�%�)aW"Y��J$)�E�D%��W"N�X%b��)�D�V%"��P"\�0%,J�*��Y	���B	
Ѫ�Q%�(�?)qX�*��P�%)�W�;%�U�%�V�+%*q@�/���_(�U�3%��ħJ|�ğ��X����P��x_�?)��*�o+�o*��+��*�/+�/*��+��*�O+�O*��+��*�_�}J<���J<�ăJ<���J�U�E�=Jܧ�n%v)�S	��J���W�{��[�JlW�.%��ĝJܡ��JܦĭJܢ��Jܤ�6%nT�%�W�:%�U�%�*q�W)q�W(q��)�%.U�%.V�"%�(q�(Ѥ��J���f%6)�Q	u���#ԱG�c�P���=B{�:�u���#ԱG�c�P���=B{�:�u���#�*��?B��:�u���#��G��P���?B��:�u���#��G��P���?B��:�u���#��G��P���?B��:�u���#��G��P���=B{�:�u��#�iG�ӎP��N;B�v�:�u�y;�h�����v���OM �ͩ���#A��:�i�?5��S��2�aZ�OZ�O��dZ���y�9��i);��SrA��1-�"����w+ �g��T�4����-Téj�*�9L�LL��fq�����4�������t:�4&S)�T�)L%L��&1Md��tS1�x��T�4�o�T��
���@�LyL��7�빙r��h�S�Fq�S�Fr�L�LÙ�1�`C�s�AL�p�,��\�S_�L�>L��z1���L�����;�Ncrr=S*S
S7&;S�?y"�+S�?y�S";������y6�hvF1Y�"9/�)�)��,L�L!���Af���Ig��)�D�V��Fq�S?3��t���ɩ�����!R)�{�T��9�ӷL�p�ל��� �����o����s��2}�E�©O9�	����1�G��!��|��OL�1��E����Lo���z��e�����ӫL�0��E^bz��/0=��ӳ\�����ӓLO0=���|�S���1=�y3=���`��i/S��é��v3�b��O�����A�L>�{��a��i�v����د�9ʝLwp��L�1��t��L71mc�����Q�g���e��i+��\�*N]�t��wG�ӥ�w	��L1ma��K^��&���c�̴ɟP	��O�:��B-�l���	P�?��8ӟ0��i=W_���2��'T�Vs�UL+�V050-gZơ�r�%L��	U�El!�\�T�t�|�y\��i.�����0Us�*�9L�LL��fq�gr�f0M�N�s�2����tn�4�����2Me��T�w�&���&������?4��t)f�ǹ@qj�Xv��7�
��A���3Ay��FP�?�4��͔�4����8�S��1e�S�F�c��������c�AC9o�`L_� .9�#;6�#�fS�ޏ�З)���a���z1�d�`J���Q�����9fsrS*�Ka��dgJf���%�m�@]��٠D��x�8�X��l�f�b�2Er�.��0&S(S�4sI;u&�I0��5z�C�ht��Ht��g蟀��?��� ? �����;��E��k�+� ��/��7�� >�
|5��:ǧ�'�������!��>�����m=��u��M��z����k��ЯX3///"����.p<�,�3�O[�;���s<i�s<a��xuC�G����u�� E.q<���@�2����{�`�����y;��̀�7b�㞈5��#�9vD�wl����#p'pp;p[D?ǭ�[��Q�&�37B� }=p���ubmE���
������]�x��Ot\>�qQ�\ǖ�����ب�;�ճ�l�ٞF�Y�=gz�{6l_�X/"����_�~���ֻcC��y�x�n_�Y�Y�Y�}��~m�jݣ<+�7xL�������� 4�l�=r�g�g���Z:yi�R�R�)��-�h�oiݷs�=��^��j+\�Y�Y�}�ga��|4p^�\O������jO��jOU�Oev�gv�LϬ�3=3��=ӷ�{ʲ���Q~Zv�ǳ��35��3e{�gR�D�D�'d{N�^��=�S�}�glv�� ��n�n�n�M6`b7���"w��m�����Dv�}�]��Nv$k�����I]Ţ�gv�����R��N�ݷ0��K]>��uS��K����hKt&�	�o�J��g8��#ѕQ� �	Z��	b��)	H���.��(��G �$�%T�Y�b�)�>���>q�/}���K�}!���S>��,�Ee��$�����[�PJn�/e�ׯoۖ�[V�k���6t�Ԅ"e���5,���O���b�����dӢ�Ettk��F㣣Q���F�����&/�V=�m�G��g�����G��ɉ���#r�
����ϝ��|���p��ly��T�h��L��˖#-��4e��q1��e��ʹ��k�_7�{7���'yƴj�R�vp6p��	l �뀵�`5�
X	� ���2`	�X, ���|`P�j���� �@0��f Ӂr���� P
L� %�d`0� ��"`0(
�| �� n �
�NF#�l`80
����  ����@�7��	d �@�t� '� R��`���@�H�x �b DV � 0��!�0�i�U4@ D�>q8���	���8|������
8 ��||����)�	�g�c�#�C��}�O�{���;���[������k���+���K������s���3���S������c���~`��0�� � p?�h� ���]�N�4>�^��n`���#p'pp;pp+pp3p��������
\\\	\\\������\\ 4����M�F��(��ֿ��X��_`����/��ֿ��X��_`����/��ֿX
`�� �=@`�� �=@`�� �=@`�� �=@`�� !�{�� ��{�� ��{�� ���_`����/��־��X�k_`��}��/���}����~���-[��`&-i�,"
����e�-�d�O˨_�h]F��{4�΁�J��v�#�h?=Co�濊���j����P��n=x�v����sRq&�1O�����|_���v�%$��V�Ux�.���+��a2�m��6j|z��{��q��P9M�4�*����:���9��i-4R�7�Z�f��C+��Ki95�
|-�^Hɼ%F��V�k��5������u��Y��5Fz���ē9��6�b��C��F<��t������T]@�9_D����!u	�.�?`>\NWЕt5�ŵt�qޫ�5t݈9#��FC���I�M�нt�1�U55.��.��C�i�b��m��}�}k
�t�g���"0���9(�Q�9�(��K���zĩ+����_����\k��:��K�J�+�&\�Ju34���C[�mF���nó��P��s;�t'��]��v��n���'�f��Nڅ'y���ky��w��6�^���y��a�y_��|���>N?J�!-Kq�Iz
;Գ�=O/�H�h\�F�ez�^������#���S��1��?��:�E��7w��͜L	����֕�?��V�� �Oi]�O���
7���iW��p�#�����5��k.�_�.�S(��	4���m��>HV�Ri�ؽ;!?��/�a�@4r�c!!���&ͺ'99ǵgh�=��E�ە���#y1��cGdY���Ƕo_��5���?8��O��Gա�=�C��-�zL�����qk�[�$)'3����2_�D���DLZ���(-44>�ս�6�gư���ֆ�pu��ߐa�G��jz���dZ��\�O:�mp�LlNM������nI��F�ۦNO�?%T�͖�^�s��t74&%!1%�b�MILH�	=�9��w樟�L�?]���2#��~u�E3����&u�sJZѴ�8�)"��h	����?�Ȧ�n2F���ud���zش�O�)��$�}/�h�|W�M��j	����ovE@D(�N�*�&�V�i\ݽD���!&�pe���=�n��H��Ej��q���]���ؔ)���rrrbG��ʚ93�ˈȘ����b 2g����vw*BF�_�>f�8I*P[�LD��KOL1�XO=M��]�32�������4S�E�����0Ӣ#�����\�Rң�E�M֮=S�}��LkŇ��S�Q&=42L�r��0k��eO4�#�,�n���rd-	�l��iNŜ6���ntJ&Ft�ML �3��;��3���wb�2��(JY�F��?n��ч�� ѿ9l&��%D������|Ӻ9-�Ed�O��h}w��Mjj}v� �b�51�ϔ�C�nv�$f���	񩚜�rxL����h�sO�z�+gf�//�[̺�a�4iɤi[����d��e%C�C�C�=��ب��=�~{�M?�;#�����-.�gVςM�׭}��1Y!1����� 2]�} �t�1wJN��K�x��0Xq���XS\�(�m��d����l5�9�ɁM~ ��0����{��h6�R����|�i�����(c����,�GQ[���!J�14fȰ�i��!/W�*���n����_u�ݻ�H����KvYtצ{��ݵt�v͝?�6���tvO��|�u��s��3�q?f
z��C���=����=�g�W=���U�@�z�h18g��Kn��1C��/g������/x�%=A�!�_le3�,E���Ub�n��'�Q�������1֒�_��=kf`uc��'�u�p���er`�Z��b6�r4D�-X;�0艚�X�Mcc�$K�=>�c9:?��-.6�zt�%�.������z)ƫ'�c�Wh\`������x��+�ۚB�)���θ��!-����%]�x[d=3�ݨ�ɢ��Q��,���(�m��pB�զ�FE/E�C�������v[��I��-��ڷ��Q]��KI3�f4z���e[��ؑ_�ߎ-ǱM���v0BB
Ҵ�Q�Z(m�m=}Z;q�νJ[��ޓ�޶Џ������@	I�����,;�B{�����=��������X��{Bp���Ӝ�"8y���zZ���G�1�`ܗ��ګ�aY�ey~�\F���#u,<c!6��SQ��E/��Q�b%�b%��>F�}����p�z�o �@7d��O�:�ux�Hf����8D` ^6ڤ2�&'O�G�mh� ��;Q��ã�*�[��sRf,	{:"%�eX�H�]�C�M<��)dg`b���(j/�aiv��[�_��Od{�}k���œ<OiK���t��[�������'�U�{������(�M�6���'w��`�ۍ_h4��Tw@d'�������fG0�(�ր���^������AV1/���U@�* d��1.[���c���9z����,\Ά�,���/���X|���� ��٪FC��9��,�"��K�)��,�~�.Q@�8�'�G�FY����`ֳ��(����LG����,��!�Fc���Ys�(8�C�k���7k�!zp� ��f5D���^:�~U::�>�.+���k[����ǳ�a��l$�S�)��c�������?}�MǍ"� �,�Q�&񒁖���+Dk��앷�x�
���t�w��"ߞE�=�r{��,��Y���8jY�
M��J��<jUÏ���x�>�D3�T{�-^�9�"�'�f����h�v�|M˻d˪�I[��@��]�>�N���lɤ�V1�BL{B�,����AT� �u�:�j�v���$�86}R��U{c#޵%�fM@���N��
�`��ϴ%�i�
'���h�b'K�ġ��.!h���4T�Ȑ�������(�I��6[<f�(�� �v�'����������C���_et
�"*��9L�h�:���?Rb1��	�O���
n��%7�x�{�Ĩ�hV̎^�ʫ���nV�nFf��jkS��)��S��))x
�yV��j�Q����4�VN�a�dX�@TZ�l*�2��V�E�!m�H>�����-��A�+�^���1�z�<��nLՋ8���n��4}f��0�T�x%�ɖ�������lq�7L]>���0�$P�@N�4|��|�z]�������0C�!4�PJ���4���9����,ԣߣ`ޣ�I�&=��=O ���� (ǂp�ƗJ���~�hGA�8�
���_*)+rD�(+8�����9�����=p�7��:yg�|��/��~qS<����zpc����g�4�Ȼ?���6���_�u��n_}�Ol���ۇ.��H_����.,�}馐Z�Z�Z��jez����!�l����X=�w��gn����0���,s�2�V*b�JSϞ���x���,�T��B����s�=���^��C��r����W���-��_���m�!���]�Z�-O@ ږ�p����s�c}S)�O�D��IYW���k�5��`�A���xs:��sp���bb������b�|2����k lca�	BF!s�h��"n�*�5�`��V�r�^߄0�G�N:^�v� ���EՕy���G�/��U�/�}������n�����x{ժ��cfM�˱v��˫�������G�����!�����gkZ�F!H�r�o_=v��ۯy���)���F�������4�4M��MQM��M��M�^��9�g<�Cۂ#^�1���W`�+6��oW-Ҙc�9<���t��GlJpA�O�l�T)�Ȇ>R��M�%��[�����43!%J֒`�j󐲹I�`���h$R��9�q����R�~I˵%�|Q��p^�:�ܐ�5��̻���5�l����������a"<��2�A~�"�+�wvuln6��닿��O�w�hu1�oY�L��9p�
�������sF�w(��P�ܡD�ŬDu.��	f<����P(J�N�u� ��8�4qB�9'�a�?�D��v��,�3B9��>�G�&�TDr�kr��y�H���&��
���*>f3@aX���Db�+p�b��I�`�z�j�M�iG丄z��n�K�_�LȠuB�z����D��|��(��ɩ�=_���9�bc@B�1���X9�J��z�h�e�=�$&�Z5E�j�f�ݓ͍k��+��b,�_y��RV_@{�n�=Mk�M�[�����i��h�
/
&��u���p���T�ml��F�� �,�@ZY�����v����#S>�k�����<S�`��VX=���ȼ�$���G�nʍ�%O-&Ƌ�C���T�����58R��AT@�𙯔Q�EûA�\�q���
Pۭ�mH5EZq@��� t��5� ���z'�Dx����5uxM�	�M�U��:��L�����	��������[FH�%&Y:�D+$főժ�U�R�+��&\��6�>ip�}�j��,~[���7$��q3�5�=.�YK�qw�j!��9\1�P����M��������3'�f��Ccd�<K������N� V�/�BX��8/ڢlD�@�9�-��3��d$쮊����v�v%���?nO�'O�Ic�8���� 9Ђ��'-�QrJ��/)�F��҂,�
��h����a���(�F)�r��B��X1�E�!?I|��j��U������T\��@�8�3�@Q�M�k���)���Jl+RA���1����X�����qD[_O�_�����J�3<N���S)y%�>�[	�Ʌ_��i:���.��P��a�by�rQ����t�ک���0�Bf<����j!�Le����~k>���8�ƺ��͊�O7�����O~��tOuD��k���u���昵�����8���߰&�!O\u�-�V�[�]	�pDĢD{N�Z�$�Y7�,�&@�[��|�u�D}���1z,=O�/FO²�1�����Q��o�'ޓ�ix�	4XVq^R����3y��Ѱj�I:rSo߁�Rrb�š	�D����kG���{V�M���j������𻄾�>��?�� ��;�~���xC��m�On�:�	z� ���(8P +���Z�@d`1�0�Z�a�yZ��$��%#� ���*�iI�m�x^�L�]uۏ�<�������v?����=wo=ti5��g�:d��|���;�5�}�~��7������u�z0�1��'�L��+�쾧����^�%�|A��"T
�_%T�}O�O��,TW��cTnͨϽ�@�h����t�r|���p� �Mɨn`mZ�9M&�QS��9�����9;������Ȃ�42Gfr1�s9U�y�F��M۶/-ǖ�e�U�%p��:#�������Z�����������`�Ż5@}�jp�i���u�W��pv�� �~�F�������.��|�Ja9lE��(�'��q�X�ӭ�cW��:|�y�̇��v(���g`HX�1��;j�[�I�[�`�#Rݎ������hp1��\M�!�4��7U��2��ʏ߶��i�#���,��d�q��%�񛞿c������u��&���Cprw��z�}�n��
�� �A��noq��M����쾛���a��+x߂����z�� ˴�����j&	B{AAE����U3lH���ǩC���X�w}f��Au?�C�E�Ϭ�K�}��o����x��\:&�\����ұ2B|�Ђ�d����4�[8 ���K���w �|�_��~0��A�)"�=
hIMDx�;��¿
����6gD�ͪr�P����JD��Q**(R/Q����U��M}����P�ZZcv���M��p�^;~��j�10,g3Z=<��|�%G��|�2�w��(�e��|��ƺ2�$�t)C�1+�#�rz��	0�k�/�A�Iqo�N%a�E��$e}�ҾQ�"PP�
�8��!hw�lzU���Sm��DG@�Y�-~ߣ֨I�\A�25�O�U\���K�wՌ�g����^�p8�K`��+�Z?���1j[��}����G$j�b�W}��.�K�X��C���qO0���m���杲T3�kWbW�5�jKM@�|N�'u55����+�k��L��s�#����)��
���Q��3.?�Tq]^oU�݇�[��-�lv��&��S���eҒ���۽&:"J�j�����b���k�=�8k��=Ȳ �jr��ϖ�}.����sď=U�(��[�#-X��vQu�O]�3L�Fr[%f�1��/A�
 �j�צ��V�Zm�Zrљ�[ǵ�W|=6�q�y�Ut����f^SL�"�S�\6�ͫ;>��`�瞬��(r����Fck׎��wP�@�Nl��7�n�`���)�L� R�߰zi<b�\��
�*Y�$�VX�4���#�,�;n��}�oh�<��}������]�����o����	�-���ݟ�ɡ_�{u��g�Zw�Ԛ�y��e�_��9{�i�cW ��Z_-ku��=xp��e|����k�f�W�KjAV�Z��J蔿U`����bC^�0u���]DD\��5_��l�$���J˪z;���[.K�t��fӫg���*U�*oӠ��S�a,�]�4���G�9`�:�d�O�&���[W��>9Q(U�vPJ��<k�Ǻ�����b�Db��̿��amj�ӞR����@��о�ח}g
7V��0��^��*�zC>���Զe��P�g~z�ƟO~���]7\�>T�aQ���u��^���_�Z;g�U���j(�i�u�e��K��."-H]	�Ֆ[�]8�dV*e`�R0��
�D����eޕ�s/^��^�`W��l�$���v9�9n�u4l+� �E�基�ν"_�	��Ku�-u���>׾:eh@F������;�(�Q�S�;һ��j������N�&ؚ��'���:�&q�c;(ۥ�0�G"7�>� �J��f�O��T�����c>�N ��z4�QrL��!#�z�j��2���j.��G%�}iz��K`'�>��E�m�������
�V��LM��֚|�7ѻ~r}_UÆ��U�]�������F��\�Xݷ~���j<:�{���tqg��n��t[�-�x[2\���ܑ�1�v#Ë� �;��a	�݉��h,ս���ˇ5#��( ��V#Ł{�9�ۮ�N���]QN����>Y�]�?�t�n4OiM~��k�O�R!�u�k��a��[�^�QÃl��Ӵ�w�(�� F�ə�� [	�.2��8�8[��y�܋����J^	�媎|���l����f _��4��M���n�F��n�@������n"fK��C�g���u��
e��}	�{ D5�����ͧ�Y@*��16��U�(b��6$�PU�x�s�PY4[^*�2�jJg�xU"K����!�7h�I<E E�5�n���=��;K>cu��ּ�_#7���䴂{o:����ފ]�V�I���ձ���������p0�k�٦���� ,�-&+��W�=	�\"'�2&E-ow�� y����rGO�J�1O !2�+�I�c^_�L�h��y�M�'�GRc�]M������*B�X�c��ϩX�2��~�c��]���w�c��k5O���Ʈ�Q"Vb,F`9]ʞN9�f�_�#��@�c�/akf"���*�=�N:D  ��LRV��,�+T���͚Qzq�f��lMe+���F��z#V����{�1ޘ�4���߱*S,�Xt�_ٓ�N j9bT3�ߵ;D��B	���V�U�zQ�_����@\v8�����68�����^���}2K�ሞu���	��]Z�;#�M3��4H���9?���3�"� hصB�f��8���H��h����	t���W,s~#1,WCA*S���a�e��YЍadpc\���q��c>3��"�+�t>D��i]�LSR�,O)�%Ș>;<k^��"2+��%%sg���	_�qK�ǀ��n�ܵ���pz��E?�A�JH���I��-�	�`�199���7ZmN�x��fѴѬ�-�p�> �Ն�2K�i�w���;���N���Xj�Upy���W�_s,5b8��H�YY�jVv[4+K!�-�5/����=�5pD��8ր74�vT-�`����F�@�K��%K�-�&��]'K[N$6Nf���)�'�9=c�l�H�� ��*a�J�>k�oH�l�K�WLV��D{�&�<D�Ɋ�/�By�;

�����Df9���5��3�w�HM��ޱ�Z�:ӶyU=�a����ڰ�3�D�qg�t���5;�D�U�Yv}�7ܻ�#?;�mX��	�����nG�-T�����l�w����ࣟ�vaUXv�6 6�����Fe!�Q�:�Y�q/�$�
|�wKC/&�Jq�C��	]N�Yt�+��
�ձȀ���g��c�!J�#l��n�E�O:���"�aN+�MU�-���l��m����\ze�.eB4o�"����ݓ�U��Q��i1�Lj���ݤ���Ƕ�>{��0���z������5��׮{�`/i�_������RRw���An��߿���6SUg����D��P]�6���c+�#��B���W��q���X�b��ҭ��ߐ�LN�4��kޜN��-�Ĝ0@���)j��pi@��v��D�*o=�l�ȱ^�k�܁ {8.	��$��<�D{9"i�d�V.�I]-�N�����뒛�Yѱ�K#�+D��0��ֵ�{n��&[3���f�7����a�)w���>�Ծ��h�z�1��G'n]�%��-[U�k�^�:�$�ڶm�~�o]��Z�O�F7���Oc�ؙ�cS���/�<�L��sy�9ߜ�˾����C���a.2�7���n� (|�lZ^מ�T�pXK����S����ۙ(H;����f�sy�%Q����%��ztV*_��#��k Ë$�iy��Ǥ�����p��K/��("����-K�d�E"��H�����7�&�?yʹ������*�&hl�X�� _�Ù��⫵�*�+�ٖ�	�ٜ��Ֆj�f�����xOc@O6�j�����^�0p�0�8��;�n��K�P�� �����P��w�Q�'�}D>�pvk��ho��]]՝�\R���^�Y�y��=د�W�.��Fr��OQlc��VB:6k?�uO#@��HxW�0�+W9
����8Qגk!�-�����c�������*���Jd�����_�{;�
W�0�y�� m�3ƽqk�Z .P�c��K��U��$�
(9^���\3�XE�p�b�4(�y��w:��A]<���������c�_K�����X|����V��k�?��1�rm����ٗ�O��Z��-+r�ǋa�"�B��j'v�����g�0	���4�#9�c�m�a��Y�Ժ';:<J�M禉����M����g�����X0��V��k��
�^T��HU���ǜ�ܩ���S�	��a���47@���?��p��^�h�J��y5C���.��{ ����Qv+�p�Oa-�ZJ)�*z��=>2v�&����[��>9�xj�{���rY4*����h��7���1�(���c���:k�:��0����2y���2, �[䜳;ѹs��v��i�!�|EϮMZ�VeM��^����k����B���Z'���To�ʑ��d���"̕�@g�j��A,~Hu�2��&�f[pƙ�J4�Egྩ�0(i20�`XR��I%@'� �T�iR	�I({@2��d�N�P�8 d-u�0�x��DOv�N����JE�rN�휄�2=Kj������"C�#�g�ȇh�e�O�=p���Ԗ{6ߚ��^�|��t}�;t�=��\o�^�9{�Ƈn}l��'��tLi���p���u�2OW=��$��@�'��dݪdc�qg#)@�(��c@���J��֭�f�F�(���݉o$� �<Ԑ�"�(E���*�
���~� u7E<M�/R8E��/E�7.7���אR�[|�J��/'dA�:z� ����>���$_�� �!a�@I�K��䒕z��,�r�G�/h���O��HnzU��5I �jߕ���k�[w=<u�}��<B^��mC{� ��p�x��a�v�^0��]��-�����{����:�õ��&���'�h؊}U���HX:�,�w�"�
p��o���_̙��-a]���)����\?
�)�'�o�2����F]Ag�E
�r.
e��k�U^�Z�%y��8DZ�-��3��3<�a�*��yXA`�INHo
�_5���Q�TZF+�G����q�� CZd��������
N�a����f���<�UU�P�ƌn�,�_"F,��V��=��5��R]	����^Oa������ߐ�s�ݕI2T)�9�Fz1}*%/��M���6���o�S�@����ԧj��l��Ò���Yڦ�H��̀ `��Ә q�4�Uk�u���5���P��厩�84�X���$N�>�,>п*�嶉�w�0�j��v��n_��bI�I��F�>Л�OZ�h��it��oe`�ߚ�T�c&�a�-��Çw>�<�Ӧ�K���Nag6�@q���?���8t`����蝝�_8��������=�,�KPu��!x9^R�Aaz)ye9�(F$2跼�F�~�{����
�ҡ�i���(,4����	^�>V��%J�� �%��0X�X��ei��cc����\�充�q���.�O;�4B�8T�
-,��R@��F����L��t {V�=��(��x	{Ei9
C�W�UwZt�tz��s��'�!�l��Ը�#�8�RF�V.�i�ged�i����t-�ݨ� �>7`���
OSO4n�!,���B�kY+�����)`�2�ZMa}�X�p!��&��xޕg+���|"}B*����k
l�.H�u&Y����E|dK�����ŷ������m��T���t��0x7�e��Tq>���6������ \�=�|�N7�M ���{<]��\U�^��u�����Y�l�����
C�m��~��.r>L_H�K��%��s����;�$�H%����l%�/��.����t��j�f�Z���S�^��k���~��d�/����o��;��U���|f��4d�ٱ���	���j@,�ζO����U���v�p�wzb������d~�������:�������*�7\� 꾐�=���]�`��f�������
����*��r�
�^N�������D�"��w������\ kWյ�� �D������Ôx1�$��:�?��P�O����.��z�'��1�<�v��di���*�����FUc$oG���\���S���>y�� "�#��C	��X]���R8�O:^H����+�
�Gpܒz��4%�i�Q�;j��lQ�'j՚>�};���!�NM��#��i&h����+{��\a�Vk���0{��S��1���\����e���FݏA�t͚��ЎsՓ��U;���O��v�����2{��*U���T߆�u�U�5��ڗ��Q�y֫R�>�t����ZRK}n��mu�O�m�vp��@�ݍmHbB ��0�d2�f���`_�d&��a�$�#BB���7�		�6a�3�y�{U%��ն�u��.��U����������UG��I���q�K2��Y��^�&��M�`[7�
���\U@��U�z��FBx���5��
�Q�W�~Sco��kUm��t�/�P҉��2di&YJ�Z��쌹7@�����k��a� ښ㵇%��x��6I���8�
�rS����j�~�&�f~guz�0T���Ih���3��-H�e;:D_����s��n�r�Z~zgU�-�CU��D��`+�u-�,���U�rF�߷�9�n��&#M�
�V�q&�ތ��~��O�qxs^��1cv3*�֒�T��w����%���,��{�Y��N��B�W!�6��Bv1*�����6v�,�������}�#&��grnr��|�L�O5��"�XwI�L���S���OU��}�>������X��v��#�l"]m�Pz6�-K�ߋ*�V�wH�m'�A�:!��!Q��(P*(
&{����L�B��r�D�ؚ���eA1�MHP�*%��.j�Vu�ע_�>�A���hn��;�Gba#c���@o+�/��@
�����@Ζ<΅�-���c���?=9ħ&��oR_!�rJ}B��Xa����kMb���*�f�T��9-ɳMˋ���F=���w�6!6���#�t�8���X�k��=1)k���I�U���v��tW\��%��_~�"��i�8y����={�x�xE�4�)���Ν��ͧ�\ς?y|�C�4�an ��Z��(1;�ߧ�?U����6����:W���Y~�d�d�g�aQ}�.�Ш�ECV/��Ņq����U5>wKU@���Ua��p�>z��.{�.r롼�=_!lj��r5���P�9Q��G^aD��+Ι(�/[P���Mk4BQ<�׵N���Y�e� 
�J�����F}ڌ�ĭ�f����1�a4�X�:reK�8'4�<-;vu����M���� ϖ'0���z��,F~�!1�����8�u��ċDk��P7�q@J�͛�s~����\np?���cg;"��\��汝����r{x�Z�'�(�P�:Y�I	H\V���o�F�L^_P;����Ԓc�����w���YVJT��TȰDSP����-&ř��)��sc�4��!�{�a�s�}y��@��c�����*�|?��z��	}��8aX��bQ-!/"6����v�\B�O�*�68}U��8$�ͤ�W7�`Ms�Ff�US�`�$����h٧WQ�RM��(��0�Gը�$`V�
��M��湨Ǧ�')4�/���v��Tv�4�H����2���R�X;/g��!ƨQF'M�F�+�_C-�<�l���\�(�u6�c�A0��5���H�R�����ȧ���С��խc�<_�)��6ƫy>8i��E/*����Q���QSU�ꩣ���֛�j�t��|�*���Ǒ��^�Vh���FŻ�P[��ݱ^�k��*�.���Ӣ\]|��rYj���$^؀�C�TY��(h)(j��f�WX>�P>���ze]�m),���ߖ4�����֖!�Q�����C�4�p�B�̙1T'0��× c�c���F�բT! �_=��*�f��%��&g�
S;աR�|6����-���ۭ��(P�ԉR�s�s^6���t�=jjWQ��?�o~�f��K�f�Oֿ�;~�+�iisQ�|YLC�;.���J!BQa�̥4���_���Տ�L��l�_P��o�|��W�������y!tQ,te��'%���w,���g��w�@�լt�ȕ+�Fh�3V/~E��x�HIGԃ��aOa���=7�����7Fg��������ۘ`>����H玻'�c~��l��g�},g�s}���7����@ҡ����=Cn�p�ٖ����6/g���YRK�mZܚ���w�z;��ɶu�b���SْѨ��7w��$������Y�/�jg&���xۇp]	��/R�@�����8�^�mDք0�2�R0$��lo�0�ѧ�]�2�0֥Ά'o�"�Č!��_��m�24]�A��2�atqI#�'i�-1E����q�U�۵lA:i����z��	!��n��e����GK7�$����r	Irl�XR��*"��lW��l3����,N�kݞ�=ɾ�i��'o<���clt �_#.�����e%���4'G�h,}z�C/5�L���RIC���3�[�O���`�����wZ�ӗ����H��Ёr�X��'Bs:38��꧋Ψ�*隕���,�Q�sT-*�y��\9��\~,gHH���6�9�F���Ȝ���0�I��D'|l���q���$�rϐK�����)��IyN�/�+�Ơg�L���jZ���j�Dg':� �I�\��բ|r���&����m�?�~�ԡ�S��P���T���r�o7a���h����i����Mw��JQPl��� ����b+q�(��"����;�f���� ��5��)�7�£���նOe+}+���a��Ax�5F�>���B-�PᾖF�BZn�jvaղ��1�xB7�M}��ֿ�5�0���HRAk���ݣ��|�����;�|�nM�Ϲ�֍�e��A>��)r��#�h�V�d�Y74vl4n�vG؁��";dڿ�/�;G"l��N�?�K��K��\{����ē�Vx���q9=|�7$�Q��A�#!�"֥��t^��(�u0[�R��I�H��O%�+rEfBm��k�D�@�p^��b���V��I|{.-�^x�-_K�LQ6�J���F(�F�ۃ9�Q��,2�M��nI���l@޴5�W���Z���	jPD\yJ��z�4��{��"�!���\C7���W~bi�����S�7��A2�%3��_��"fW^*'�#~��;.'�?CƉ����6F44\\&C &���щ��\����\�p�cp�\�U���C�m>�!�~͠�ugc�龕�	lQKu���>`h=)�:ZO�ȶR�Fl��;��έ�:�mlY��<��{3��g��~�Y���mF��x�Ɣ�c@��YP^�3/")6�����'�|B��Dld�������f��oD(��V���ͮ���6tX�<=1�U���C�Lo%3�l��fp�>	�F�V"�:����S��8#L��֌���dq�� �䊬�ؤU����/�.
��m�پC�B��pm#پ�u��ap^F5��J���v&�ib,�����Ễ�V�.�?i��wl�q��є:5����^ .`��D���\��5v@��|:��=B�ބ��>/9����f�S�HEf���^���+q�}JtuB�5b���XN��]�:�OL]�5\FLH�]�3D��~	��PG��t�� aI� �15��@
��@\~�%�2
n|9-�6A9�C9?Mj��y1���D����� )U͢�iYsu��y��{��q{B֫b����e��o�v���;�C��o�C{g`(t���{G���''��u�6�>���sc_��{��﹡�s�D��jǩCꡕ��䕒�n�$kZIִ��J���0�&.���%1F��^��*�
3��*�+/��W^m�d�[{��C���R�I��6�Y���ڔA��k���$��я�m�q�����{ǘPg�6$[m�o���é��m�'�l�{���v���ynp��8~>��gD��e�����HM�Z�����4Z��":DA��C����vH��k2lъn]گ`��>��^�&��B�K�5��:W�޺ƙ^�$_�lIF���cl�t�UU/�.�tlg��a,�����
�kgdʂKɾ�I^��<��wqq�X�Z��ɯ���b��b��$�ml3"��I�k_��� 	$ǄJu��I��L�@�6IHCv}ҍx�T��g:�Qj��V�����Ԩ�vo��l��������>�!���n�|�F�Q[��=�\m����(�V�1"<�M����&��~cn�813�''�&��������廖������q�13[	�-�@���4������v+�a�W�?�'���Ѿ�ndw��,%�-�a"�s����,�,ϣ�D�`����R�'�O�}C X��������q��i�u�T�A��ږ���L�бp�t���V�p����zS�w��q�R<9{t6��'m*�����J.UJ��٭�Kq`� @)�;��:�����:�Pz���*mz��ћ8�WrN�n�Ļ�Pjp!r��O$"� �j��_{�����"x�L$i9�	�������{�-&�ex�b�nb�(�)���[�xcv����Y*;�����|l�����S�0U���(�ш�V��?M���d�K��L�Y,�g~��Dp�Σ�Uo4;93��f!g��v</�����.��9MU��k���F�L���׼(��j?r%�lW�oӚ�5�����B��'p��w�dF8�qf�'#�W��8M�k���W���}Cδ����w��[R�B��r�HJ ��ә�@�j�|9Y�|-���ʲ�Æ�R��c�nZ���@H;�#�+�I�b��$�pF�	�Vd$[����dW38�g7d�a�k���|#eT��g����E�46]����P�*ߜJ��K�eؽ�R<kp�ܯfɬ����K��G���(���3f�x�jZC/O����B��H�g�C�n�8��f���;P�ӞX�(���anz7����MW������Sm���*�$���PzR梔=�$�p�i3����tU���V�،��
�1�B�2��i�]�p�F����he"S�a~%4�֢�4g�g��s�� W�tY��u��T��̺5�5'9��LBȥ�+���_'BEFɿF���%zX��8�fP�����&d%�TWz�g�Ձ.��<�҈�X/A�r���Jb��]�0P��V�$�󱓄+�q�V��4�N��8yqz-w��t��r���K��*~
���Jt1B��NO��:e�z��]�-�4?��v����joF���Ѥ�H�/΋���(u__#.��)6C�O�(�kΈ	�h�ȨڱL��H3hj��/�jj+�6`y�VvB�C5+f⋾�p�IJe�%Z���<a�W������g����V�z3X+k0�b �f�˭�j�7�%^���������q�|[d=�B,���mZ��X��M4q���Gܪ�>0v7�����"$��)TF|vp���U�_A�
A�!�$��M)}��.��ڪPo�օ�p+?7�Y975��?'H7q�bJ�(�K_���֪s�
���z�_�KAk�*���M���栘�ok⦊�[H��	^U6�K�" :2\}��J{���,<جⴿd���E<#ZD��-�rj�^q��h½��ƽ��{��{Ua�ϣy��Q�f4��wO�C|�O���d��Fy26�U�@Q���2���ʸ7�m�L/4��"�
Qަ�V�&{�P��y�ܿ��4����aq,&G�v\����sMb�0*Tv�*�+1qm��\��x�<P߮����@GQYEeq��QO&�<��xN�o��'�<9��6���ȕ��!�_���x��%S��hg%r���X
�^j��u�4���Xh@<�@Ү#<�H�u72s�Uf���e�S��A9�f���CG7��~�l��g��:=x˃7��z������m%�4���]�uR�$���o��h�ݏwr���O��8�6��ژv����~P�_�A�I� Ƃ84%��B A�g1"A��@$ �&p{<����� �����%t��W!~Q�zxa0Q	�\ݤ��iO����bZ�������L�}���7����q�P�$㬪o]�4�## �H�( )�v	cE�N�����F{�ٽa�FQSP&�����cUԗ�^�����!j��ڦ7k((�$|Ѽ����_!�CR�C|��'�>ȗ /�e��wK� zQ)R����hĂ  1?��@���P�$��@?Ȁ�6�l`��� �{Iş	���1z/��t��4\��!��� �1F����tT���Ϸ�6�]��`,K�m���}��?F4��X,^�49��,��O}������?�n�Ћ�)�ml���$���F�PT�m �~��r�;ѝ���0/��)묓q,E��\l���OA�ޢ��ϟr��䓔�������Gh۠�	A����_��u�oV�?!�ˤ�t9���*���g�3�;�\7YUd�� ���@���8���C>"�Z(I��Pr�WD	�C*��Y�,�iY���p�+:�]�^��4HSR(w��$@ot�.��#��:]�=Y	�Xo���@�����)bRQw �tͧ/��������M��#jK���t���D���<�(4�Q{K,�7l�*.��в~�7j&5�?�-z�B�{j�#x_Zo1���kF�AA)���)0�D{ꬦ��k��ԝ8��$R�)хl�$���Ӊ3vɸ��4]�8{Y��_qj-�b����xhW��hN�YA�z�'I�9D� %R��C���ux]��ͪ";>��\�Tީa��߫����jh ���l(�����Y���V#�S�����HSj��,��EG�1Y��A��:O�El�o�)�v����r�Nͨ��D��|�ɛ�8-3Q��-&d���rV���q13�.F}$��ڨ~�e�I<�L�c��K*t�^�>�_U�x��@E=�����7E��J#����y�Q�&Hb�|�,�n"C��}6������*�/��%�)�H �dA{��%�Y����R�����!i�o��b���һh �� /�ڎ	D���>K�)x}����X��<,�6�<������&�&�gcr���,�}AWt��m�۟�F����`Ƨ6���׍���>9���mm��/z���Mrm�TvC��S��Ɔ=�����}\��x<�� ����1��؁i���?��� �T�%,~���dhɹ�x��}XN@��I��(�P�IA<��8%�3�tS�
x����(�*)j�M�>����8�!�3�J�e�������^�g�B$Z�%ƒ႟��*/mLk��cPo@����F����|&�۸w4:�Hv'��w� �]�s�$ډYig���c��v���i�z�-�E�a�wP���*q^�	�k
}A0-�Q�	m����eh���m�W�l�=&�B���'?���uȚN��:%�̓J�(�&'���1�J#�N�٠u��̡��RǲZ�٨�����}�����5,Z���^}D�B;�%b��8��s0�ɀK����P���R�q}����(�27�I\��-���f��[�e���Ơ�d9�2w�����\����lBe�U>�KD`t��b�J��W��ù|n惃�C3�Xdi���c"]ۜ�:GrW0݅�c����G�,q'�I�¨��3n�u�.�m%;�75�c��H>X�<�8,�ʵ$mI!�]!�����F��j� n
^H>$��G���6]H������~q�eB���"�,�c���|�Xj�jc(��	<�H||�hB�+6��;#RA���u)Ng�[\�Q��z��4�J����=��C6=B~<����ux�l&��0WbS������܉�A�!�A<Q��Y�(.8�����B'��3�DDsJ�>7ʵZG��XK �&JJ���h��h�ݡ4��6��i�O���x���ih��G�YK����:jE�z�?�����3��Rk�+A)���� 1I\O�J��l�D�0�Y8�m �����'�^wl>�"��1s[�u�DTq��`b��m�����LY���>P:ֽ��+@ �u|�v����.�2������>	���_ dO��5�^��)���M����[���1��U|���1��T ��9p !!��[�����}u,�+��w�*�����%�J�tD�1h&����u]�^��<����+'���}mqO �✡�m���N���w�m����݆lW���cb4�6)~��,iG�/�z��1;H%i���#�^.�H�9Wx����s|�[I;����z���N�����H�;΅&G ��F~���H�]>�0#zg�av��Rh��}H.��k�N��6������}��:W��&�΄����0����G)�B���o*p�֥���ej�����O*��-�POI�ϸ�$J/~;G�."p�'������?�@�uNp��W�;��\XV={OS���&�M~b��DB��`(�l<3�P��$	_Χ|�d��#��?o=|���R�~v:�'�0b����\̻h}���O�����]@��+yi�c��Zz�F�[�-v�~p@�3|7������J���F#*�ۂ:��r�p6$�o���)U*����)������z#J�P�:��/�:">�v7��`��B/Q.�=�P%�g?+˕$V�.g������ZͺkC���F����q�*���<����J�:�К]��Fc���u�&������`�^Qj���j>Y{�l{L�����}�-��J�p�/����a�s5��qoIS���q�L�������� ��C���k�O/N�-v'��C�&�Ju�����D`�0��᥾�)a�+*���+��D�et\}m�oaǰ4uvFJ��bs�T������;�a{a!_��pw�r���umU_yL:�����lO�s�"�f{%I<
��&�av�Hx�'�K{`Q&�XY��&�1n<)4��TGxj4z�,�Q�P�jwox,!�:�:f�ˬYu���.��@K��\O��X��%��j��ʠ���:5-�� FM{����B��A�^��M>�����Y���G��T��1E�eS�V�>��zkdq6��?6rpS[rb%1���t���ʝ���x��|Z��(��k�m8ʱ6�h�s~�^d��T�Umt81�i��렳�{����΋ձNqa��-���H9&��a���D9�@����LZc�Zk��h+%���H=!���}8�Iw~'�E��
`�?"�G����1*ȁJ��'�UË�����Ǎ��#b`Pą������s�N
�%c��>W������+��8�jep ��s]����!g�-�Q�86�Ã�Q�^��>5�G~"	��<>��~���x�G�E�PX�wi/ƗB&�o�v�Q���E���^�_C���n�����0���:8|��7�5[G*���
F#?bF��u�������6�O��
�҈��YO>��E��[D�r6�h�;/��%/�O{5��<��~��GG��Ǿ˾Ȓ,�}�yǱ��[�����1A�<:�����e��p���,�=$I�r�7�o]���Y?T,�z!E������@֯WR�J��&�����P���m*�:�.���\$�/��c����H��8t&��n3X�4c6�➠ݞ(u�ӜFo��oX=m`I�/��x��0�ד�DA���"��8�:c1���'������T����!.���q�o���ONKɢ;!X�ҏI!>.��q�px�2�Y!�`}�Tj9_дk˴N��O)�����H��@�S*�4I1�:=� �����jZ��/ű���L
�����]��h�͚���^4��a�\�/N�C�����W�	��ɦ���,�훒Lܲy�3l���=����V'����Iy���<t�I�������*��c�'?��Y���o�9��X�� �,>Pҩ����h8D,�C$p�\���-�/�t��Y}*[>�O��n��R<Mi�!�'l�R�д��X9�YI=DR�j�M[���7jF5B/P������^M��7;-��J��`?��P��c��^'�\Κ��)�V�U�Z��ZD3���ڽ�[g�܉E�!�gⶮ�-��e�fh?3�Õ�5�ﺲ�����'uI��
��]�MC �JcEGV-����uY�VE~�$o*�i�9�J��$yP�"�t&c������D32�:��z��( jem^'!�M@oi+�a�8$z!p�p8Zk��C�u���p��N{���a �K.�u�w��;Q���6	I=f�}��M�	�Ix\%�&:{,�D6��ҫT�F0��gQ��(����+�(��_��p9���:|�R��6��D*�L��ѫ$T���9\��5�~�T���;��R4F� �"o��{���Sj��~<x6�4���w&�mT碟3��6Zf��eٲdٖlK^4��xK��Nb;�ĉ%�
�%$@(k�ek�m/�P(K	���A�+����J	�p�.?h��A��-��l�s�F��84���^�h�љ��,��?����d��Bn�����{e��+p\��_V���J�]��UUԒ�%oǶ�T��hWQ���rXLp�"����sv�ɡ4�V2"�R~�4�u
)Q0�Hp�D��e	��^�Up\w�ӳ�!<�3�����������PQ=�.�ȌW����Ұ�} �@1�<���@��w�� �0��X���=�vM����&�����7��T�SJz�\�f�i���{�Ѭ���O�JbH�:�WQ3������wZ,�P��_��N�N�(�S������?;�=�E��'E�%��нE.�A_~�+񽷭���Kܻ�$^]�W���U���jx��>o�[ �8�.�v�(��;(-�Y����a�W���/.)]����p���4H�^�ի��d��Yd��LENg�,�r��g-���Ӹ;hek����ʮO��� �0J���oѷל�X�EEt�xF��e��:��9e�Y��Ț(�����W�y�iP�	P�a���W��,���ͦ�E|�+�.�IG���X�8iEΉ/���B4�ro��2Gn(<�%���@I�14�-.~,����%�T$��{Ƣ���V��@��.�4�o����V#�.��ZIQ�py|��ov��x3��Z�ES���jVV"I|��!8)��\���r�"�d�,��6�$`=�/�fcg�Iފ�)�����K5�}(�VV8��g�z������F����}��](�B.(X9M3j�g.{��aL�v{�,���^��"Eۈj�3�)�G���Pm���g�F��eH�%�~?�~?jx�+�Ŭ��ju���6'�������4mx8-\��/~W���)������K��x�6'Ckw�4ԁV��';�7#+M�V,���ho�_
�@DR4[Ѷ!2t�Ph�S���n�`������*h��]*>��-�����ou[ ����&	)�U����l��g�[Y��(��8@���v�M��F�o��-���`9/�cs_�J�ؤ�����Vj�Z�(���g1���]�h8d~�r�)�G�.dr��{n�����,��߫ːל�;��NZ%���yֆ�:ǫ�X��W��s+�ٝH��H�\��@Y��r�J� (qyB����'ਰ(�������k�!���(�,<V��d�$��U���:��e7h\�{J�k������p3���Y1u����m��K����}��m��(�^�(p|�h���4b�ƅ�������&)�������?�L�Nx����)�A�Ev�Sz's�H��TFc�A�MI���p�1.n�����b����!��f�E��*{�m�xo�Hl0�X������~2?�#�����~�ξ}o���"��˱ֿ>����ƬL�d��4��t<��T�6?D(�E�}�`�����Ȩ6sq"��X�\�1���V�SI)��Ů��-[D$k3�m���q�4�{积M�R1I3��e��O���P���ӊE�����iA^��5�Z�Y�!&,��~���J�P�?��.���|o*ͯOݪ�����m"�ä1k�$2�©b�4��j�������'�-��4���O���|��'��Y2E�Q�����=���<[�Np݌^M<Gj��ͨ-r�x�������ҿSy
<k,I���6�C	D�mk:E��n�s)Y�
���ó'���>�#`��I��a�JNS"��O>s���"�#{�b3|5|�k��z�cI�vj�|�>��!V+�N�<������/_�!9���3=y��5j4&��(׹�&�N濴�\�Oݼ�<��~�/[~�e��,|(��*�T[��:�Y5᫜0Ìz�E��e�M��p:�Fˑ3i���.G�j�y��箨B�c�+�f|�W�uX�u^��up]���~髃���t(��w�t�����kwݽa�����d�X���p��bYgd2�e��L�fmC��ɹ�HS��U�6���4� �Dv�/��Ū�r�Y�2\z���6.�"{�S#1˰�b�Ԧ{��93����I�X Ʉq8�n��[O��b9y�� ��y�i��[3 �˪9%��H�oơG��u}���4�"�/aҹk�袙4�
�"!ojV��HB�1��VS�80I�7�����esq�A%��J�o�К�:*귵G1D:��r5���o*�4���d�T-��h���s��.�V�����fw!��
]b(EUV��<�������-?�e� 陟���$���O��+��ݩ@ww E��r����i�L�`�������6e��=�]Z�a��.C�h�,�S`L~��|�2��	/��ht�uǄ՟�Aa��2��[�d�6���;(�p��'��l�V��/��1������&OI��Ϋj�������ɶBK�;V3�^.�37)��k�w'o���=}�Gzn�Ykp:��aК�b�����ܘ�@d�kͬ؛�TY�V��yi�jP8���k�?�R7�[� ���=p�{�r��(&u<�f3��t�HD�2$}�d�Cakaϰ�壢̈́�L%���U�YT�lZ(j��
	��^��>��s9]8�^��k5�HQж[+��0����u��[�P��6��$�C��VO�[h�aZ���;�Q��X�A��SHղ���R��g��Ԕ�G`:�ê�O���
k�l�!� f	�2jfJK�J��3�J��gҰx	*:]2H�;Q.2�`�����o�v�V��<5�|�ww�'zb:9������'w�y:�p���6��N:d*��i�k�k|�ߚ�8����j�ޤ+t�fVf�]M�m����Y
H��jmZ_`�>U9v��G�L�紋('Z�Xz�eȦ�
�EQ�!����Bu5�_wF�)���X��\䐬(X�L�Nk7Ѩ��JXZ�QŊD��	r�+~��ؾ�k7'���t��G�v6�rR V����ڊ-7)Kj�����C�Ϙ�S��I���F���o\�hO��Ȗ�'����2���Clb�*V�u�;�j�I�~�h�Hʫ4:5G��
�uo�Ƙ˩#��8��ܮ�;g�b#�!�g	#�e@�e��9j�p*�=mA��N�q��e!�8�7;�݀:�B��2��䵺�,����'SÙ����Jψ��4v�E��y$6$(��]��i
�ʾ�������L���.ä�����j/�@�+�#�����&^!����s�M�s�����/|��.հ�98�6o���6�B�WeIpQB)�}�H�++��}sy-+����?:���}uE]�[j7���_��ks�ݰ��uoG���v��7�m��6�hN�&�_:~�͠����PQ�U��&:<������++J{v�W��_������c�����⎊�s�w��nW]��dlj
��a(2P�D��� {(=]g�y�GR�@	R5�S�|� D������B� � �ɰĄ��dle��	U��d��S]Y�5O�-�n*��Eb�T��1"-����Fӏ8��xधq�o�Rk3'�R�w�W��z���Z9��ڭ���jَ#���eb⎞��_�2���=�.����k,�֩5�'���	�16c&4f�и*sLh�BLH�T���c�o+����o/z�T7�Ӿ��n��G�IL��EĄ���ƯL'S�l�p�>��"��z�#����j��1��0i5ޡ"82u9�z�ani5�
��2K@ey��J��p���x)��X���K�XP-cG�Ic����JU2�	�Ç�[��p2�?1D9ǈ��A�g��8�E��7�:l�D֟�Hr��R/�!b��i�P*���-fcy)�<���Q�3iXT[���{�-�F�J�`6~���j.�ҫ%�\� ���2vlk�֎r%��h�!9x ����s����(���Ș�n�u�n)g�Z����H���O	����u�1G�ed;�\��_��׮��
��)H�5\g�Ĵ��W��r�mÆ˦E|u[e��\%i|���R�X��w�|bWþ�	�TL���X�tSj[�'�w��X_1���è�%�:��h�EKT��o��8X�8��i�Uz�C����>������WTnZE���hM��AQm5pF�B��Y�@Q�مd�j��Hq�)RAR���
�a4�E���.�Xq9�{�x&�-	c��D�?t���Z7ޱy�N�P��H�
9���n�0������F��bRR�^m$���EN������^Ήh����hM�ρ��H@�����Y<��EgҞT���������&�%������ҵ��1�ӥ�D^�:��qoO���ځ��~�uh����۽m��G��3;�9�ИMJ%g�4VNjv������#I�b94�dl�6�vA��}Ȍ�k��u�yި&�F�A�PL$AcD�������6�������H�@0��j<�� .X�hi�:�@��Q Ef�^�(���h�E ��F0�y�x�fQ�[9Z�Ur$����k�9$m�$_�~*�}=�����+�S�ɗ��H��@{[P��������O+!��7C(MnI�[�����/�R��Q��*���������:�I��{z2��+m+�'aO�/�R=������ *5�J�&�R��R�JOb(�j����s��v��"�.���)E����,��*�+�*ѲatV�����gb�3�ܙh�Nn�-%9kC�S���@$W&�[��'6�d ��ul#�����.�i C�xbcX�(UzA�\��T�5�z;��
'х�ϒ����,�K���Y�pd�c6O��x�Zm(G�HE�MS��N�:%<t
N����cut"z�2DVQ��]����
ؼ<yh<A�yx;s�|��\`��$�l�Gwm��=�@Ǟ��aH�[1ɗ�%M���?�W���Ӑ�k���=�;��#u��7�t��q0\�{U���=ÕMWn�,�'Y�e}���HqSČh�6���V������4�ʦ^(��4ߔ��-����H|CY�ˊy���|���KX�dw1�D�v��E��^�̫v1�/]����"=�<�>U��B>�ʋ�=ec�o,!c�����TX>������B�'5�l�������X^Y�d��u:���ըۯ���3R��ށ��N�n�f��H�m������@Z}�o�$�*L�U��U3�	��S��ń���?�_��������OL�~8K�}b/:>hO4mo���נ#i:��Ά�~tǱW���oz�ރ�$���Ǣ���Q�̅O�ۢB�M$���Y7��6�ڶ�;���E$�P+�(�ѷ�t�dދ��������r��dt����+hJ$����������Yg��=&'�v#g���Ȳ>���!�E�D-1����%��9�o�l�A�@���)񎬹7~iso����W co���_��[���^|H�R:w�J��r�����:c�1\�>���¤H�U��\�[di88�x[õp�L�Q�0��5Mv�=5%&��"�l:��S����c[<�����U�V���V�����W_��<oȁ�� ����{��l�|b������{�'h��r�s9���2�$��Umi+SC��`����ĦZ��i�e?�؉�Ji:�!���J+66�P�6T�l�еW�9b���є���7�-(ٕ�e�f)M���f�ʬӘU�%�\�*2Y<Ze֪��R�鼍�����!9E�6�Q�_��:.�A@�V݈[��i�(̀�y���� 
�YV��.߉C�K5q���`�g!�G.��re!���h}>�;H���5�oHtNʎ2_��4�ׂ[�:g��	;�߀�I<� 9�U0jܞws��Ҭݤ���*��QɳI ���f�{�W����@� 	��{��G�=�e��`yEI���S�l3���K�:��M���O�KhӲ~�Eq1��/6�1�	�0L��4��b���xwEj�w�q�%�u�F��~���d
��>��b�����2�N�p-kTI8�^�h����f�bC�V6�;@\���=��vBiT�b:k��P����x-��� ��N'ﻠ��?D��A�
S�1\�AZ(��]Hk'h��E- \s��^�2��Y����}}	/�[&�q4$���˥rwY�x�t���W5�n�����������Q���-7���7�T���{ono��{�"F͚M(@W��'Ǝ4)����`��gPm=���ԬE��t�J�����CD�A�;k���\���g��ч�ut9Q�Pz��C"��kvr4����Ӱ�	Z@�\c3�}�A~�P�~��r�����$lKD�ġ��7B���K�Yx��#�P��Hd��T],��7��o
��[��̫˕6�L�'��7�v�R�K�z�?����������#N~��94|���M��h_��F���G��Ⱥ��.s�`*�_�m��qSL����@A�hm�{�4���������pu�=Uc�ն��Ov��NGyI�944����"{U4jsU���~��d'��(ђ��w�	g����I4*4Ez�%�Q8���'	OX.HVJ�<��'>J�R�qq��BZ������Ϳy��M?ݩ*l��g[���B�XL�$rZ�wE:v����T[���}����-�}���xwy�+j�����n<�1�`YF��(��H�)�F��*�P�lYs�x�Y�a�-��_��zk�7O��XGݰ���:B�����Jح\���)�������C^�Y/��	�௫���d��x�ީ�=���\�н�v��`�w-�=���R�5�S��	s�暗O��S���\����o��mק�� ����}p$�	J	��0�.g�՜spab�p�˟�n/�>x����
��^T���a1��"a�	,Z+.i�-�e�x�Y�A�1�/���
�a@J�����Ј ��6h�j�Dm�h̬���P;��A��S"
-�|v *��b;�VQ�b��25y*yJL�&C�9�W�b.�Y���?|A�<���?�_��Y;]Z�>&Ӻ�&�V2�dX��]&׊5�'���R?�!�C���~M�HD"�����tv�AA�3\V�M�Ȏ�7���P�ί�:�8ZE:�:��X����x��6�GO�Y��/�/�M]��_ͧ���`���~`�v���A��"��=�C��)�#5��YV�Ej�D��G�V.�Ö���#�~��P�J��)8�NmPJtP�E{�K["f��2�@�}�U#��=I����0&�]��q��SA������>��	E���0��j�rJ�"m�W��=���5�K��2�g�W�-��Ж�F���V��la��c�U~���sH$�Xk��=�.��恡k:]��B�����=���e�mG�M�����WHjF��*���Q2��k�ť���mQ[�y��^_Am��[�(iX���on��͍�ZV�򖬖�|�����6�/C���P�{
Y1xdeE������/*�'�DP�r�U�U��ۯ���(#r��,�[OnS:m�#-���H�%)����V���T�Ɖ�[��������7��	*�V�Z��ū*z���t�^���;F˝���+�c�������N�ߒt�4�e�>�Q90�V��:�LSӻ����Wܩm����:�)��YR�uM��i86p<b�mZ~�����A�|^G,���OGO�����>����n��Qu���
S�{<��J&LH�;��oą��I��]���K&$�r
�򝷢���z��y׽�Em5~VF�8��(�ٿ�t�d{���]���/���]_�Q}�
�zm�^[�Q�2M�S��pp�\�b�f�ά��D�;ڌ 6��@K�1<�o*�
5wA��@��������n��D{����R�M�d�!�d�|F�烇S􀠿_x7ߢF��N��P�|&\ʾ��8�/y���]{��#߻�:x�)^w�}�U�����p�����S#�_��W/�x��C�/������c.��6n�";N�$�ˌ�`l�t?Z�q��|u
��'�Z�H8�B&j��������@��s�|�f�kr���%���sWϚw�ؼӇ�;�S���杕��sً��',y���'0��W�yVs�j/#�yg�sA}�l���lp֔]S*�ߙ&�2.1��~˝�Æ֛v�'K���]c��$�às�J ����`�+�����]�2r*��g�_�\퉧��%��IP�a-�yi�Y{����Ym���-/�K�d���f�>�e;�?��s8���}{7�9)M)UL�{OK.��p�K;��7�^�,?�؆醡[���T�m;jt�J�s�V��x>���o�B�|�"7Z>�4j���Z��`k�dO�!����x�OD"Z��ob���9��tր=������_g�^Z�g�y�W���������4/Ku�[+��`1��eZ�;�eN��Z-����c��/����n1k7j�6+G~$Uʲ�}?s�o�u�l�VA�"g�ya��m?%�,\�gu=��]�(��Q@�3F��]ޟ�0��,@8�/9��T�ݡT���~N��t�P�xx���q�hdZ��5�R���i�j��R��@?��%�`���$	@l�8W"�H1�<!�M���zˣ�~��b���(4k�a�W� �� ��?$�M��n5�>}U�J)�9eZ���G.D��BL|��N8f�wTJ�ՏW�`��_J�?!���JvJ����8��K���	+�>�Ƒͤ%�5���-�پ��cG-��5v��ʊq��cì�h�ދc�~����dc�j�}K1Z�&�D0�&�+61+�mbB�a��4�'C{��Phrg�L�����g��p	�V����KH��A+�|(o�erl��ж_�^Q*_''	��X���.��W���P�5� y�2�b�%J�ʾ�99����	͚����)��Dy�"�^*��̱��F����QY��]���:��a������IF�v�ǧ�6<~�{/��Sc\�_e��{���ф�q���D.��J(p+�|��x��g>3@IT����啍���Q�D �*�(vJ)��Hȿ]$Ty����(IH�0��Lze8�����	���ϣ[���2x�C��)$9��-b3@��d�@����[w�Mp /�#ޜ3�$Ϥ�-��K�����*G��>y6T�E�&��z
�"�0����DYT	�PdG��L.d�4اop��dh�-���`�UȠ|��-�1���˹�qf���з"$���q�-��k+S KIKM5�v�d�����d��C_�#�8�j����&}��ur?�>l����Qh��AX�6Tу�L
����2\�e��ˠ���ך���G�������^$E)��5_iEWZ�� 12t'n&��P���n�F�
5�6��mX[�ㄿ5 axd#2� ��t�8c����MѶ���R�J Uꋢ�R���/1��X�M�O��1�`���&��v�
�\�V�˫6�y���*�V�pP�N�����hU�F�H ���U����	��=
K�������V����
��o ~=�� ��I|4��@�
�,�dei�`��\���{v�_�C����a6��o�%X4�YԧX��� ���ϑQH���T�"�~,EJ?����Aa�`9Wq�F��?�Xئ��F겛-��V�*i����9�(9�s����鉝&��w'ǝ�0�9i��V�jWBB4H!!�d���p���9~��L��,`�Y���������]�g]���E�W��3;�
�W;�5�3��᫪����9��<g�}���vj�6�!�z8��'x�������y���ޑg��!j��>���`��d���S���Լ�7�ȣI�*�4�iRֆ����=�C)"eGaGa�ێ���4Hc�	5��L��P�T���@��^�����;�`�����p���t�ox�.��a@����l/sUO�*�r*~�y�_L�q����3s�?⟉������șZ�Yx9h�-��M��/9hB�,yhB��C�o��vL����u2u��s��[��HJP���>��U���bz
v�q���#�w��]��j��z��\J~�np�oq�{Ct�3H�� %�0H�	_�>��\MC�D�6)[E#i��>��3��X�sl$U���ڸ03a���$�f:�43��!���w�J3�ߋ������\� P��HY�I��I�6����$ޑI^�$ڒ84�pΊѴC��"���B�PB��ZBx�G�__�s�����+�9�V��~�_~��rDФH!M��UO�i�$��7�j����q���x����8]R4�K�\���[���ֶ�ҮW"�7u�ke���x�xz걯ݵ��fy�i1Zh��t�ř(m�̪��ݲ����(�a0~M�P2"ï�/x���-��K5c�U�ClCI5x�:�F!�����4��QJ5���kX��jfa͗Ż�RM
޵Il�i��<x@l��j�a����j6�Q|��jX�K5Ӱf�X�C5�0~�E/�fDʓbD�("�K��K���E�|�� �/U�G�i���iӢ�]����[֬�i2Z�^��`����":k��-���{�����o��}Ws;�۶jO�=8��_m��b��s	�z0�8���Ə�v�p�I��M҉���tb[w�*~�<�M^�{�zoE���h^�v��	5D�z�V6G)I�n��;I:�U�{p�ѹ~�ñs9��4W_9
R��Qwԍ��@oY�4�:�ɼD�X?\�X�i��ި��KUؠ>�+_�w��4F�CC�"j��Ъ�����%)�RȔrB�GJá���Nml�ȕ������i�k�q������r�����@�
Q���������5��N4|�������`�78�+�y�ϲ�G#e�e8r짎��� /V�#1�hh�:.��guD�U1� F�VI�X� ��i2�dS;87�[
qs-^UM|+G��k[~�`|<�B+�*�ܕ����Éa�
-"���Uӝ]���N)Aj�KÁ�]��e����P��ti8�R3&�h��\g�w�r�r�yo)�әt�]�k����e�چ����'�P���4�_��?�Xw���%dw��K�l��jK�% ��;C��i�v���@^{�8(��Ñ��m!�f����|���b�R#�d���A��S���2�¿R�9 �L����7N�nx�ᯖ��<��P��/���"Koꊞ����h��jt?)���m����YLEW]7�d��@��)s�'��}�P:����Έ_q������ń���dys�WAs*�"C�N1<�xr!W�I+x#�̤W�&��:pgi5��_�����U������O�A�Ï�M�
˰�n��DH�܁��[���%����*l�y^�r���/B����}��:��o�:<��l�82˯3�#.��<�ٗ����5S��i��ve�e�/�f=L,�q(����Ķ�WW��B�18��T((emRo���uy�^���ə��4���M�3����(���u�9��c��e������e%a�_��]�oNBl`A(d��	��a������j�J��	�6�hϫ���B)�J_� {�6����$�΅�p�X;։�[� �8�b.��ʢ�[XX�g��Є���e��-E`^������������c�נ�/zb�l�>V5 ��U��6��Iyo���[�v��_��w�Xhݴ?�{�w��o�q�����HwO��q��{ͺ`Wȟ��#��G�]W��C[�\8^p��e��@��r_�r�/֞�.[�=kz=:��4e�q����ZG ����8M9�Ǖ���1Ȕ�ep�����C�/���3z����S>Z? �B�� %<_���sْ�����1�5D��33�g̑��!Xj��.��+2�D����;����H,�z���zڝ	���*�}��O��U*������&��
oem:�i(\��be�`6�6wƫC�7Վ�[�/�P���b��O�xI��'N��g~!`�	T!����N�,�0��&m*;2\-�ެ��}7�К8ެ!���>����>�f�@Fʺ������C= �8������[/�.ӈ�tP����K��IƢ�wL��	TS�!bR&�CF�5b�zޛ�J�H5Q��(�t���㞬O�����=h1�ƿ���}(=%4�����#��
�����h���1��5��c�!'��c䭐��PA�y�%�z��"�Ǫ�ÿ��	���5<������5�|W��֝�{3nV�#�vj�eץbko��y&���q���h�V�g�Gi�h�܇�m���h�XY%�Տl��Ë�jY���GU�K�j"���Հ|!�*á~F��X��!9���������*�n�8d �T;��Z =s�T���B�QUeeVɚpӱ�!���c�'mS"q[#�B�z�
�cUئ�Y��f�hU�-�R�o���\̓Z�܉$H:��x!e�\x$���ڬ�1��1���Fo&�n�X�]�^��y�5�v��-�N��5
y��Ϻ�\��,k�������a_�@�Qva�l6�&��#}�0~��0z���;����G%�1U�=s�����4	����#Ug��j�H�����#��K���oa�bX64���ӓ�3r�Ra�tF�I'���{)U=4zeh4�aτ�r�8A�|��@aeު������hƮ�9�l��G�f7g�Y�(7�S��Qo��12��V3�J�i�m]~{*lW�,!�'Z�C�����,{G�*�Ơ��c�H�������~��T[���xVׂg	�g�4�1)5U�?�= �Q�?��+؂f՘J�G���Yl� _Z��N��gU��2�<��ׄ�~����=���
u�藺$~贯�׮��A�0����䅅�q4|�ӈi�'d�Y�l����}8~���4>��W��Xl��p�.<vE9R�٠ �r�)P�:3��H���1:=>��j4����l熊��̪�S�ժLĳr��Z#�TF��q���v�]8nNc��{ 
%
����?�&.*�Q�QH�C!�uᮇ��.��o]�M+J<X���CHg�u4W�.�f�`6����ٿ����qV��k�+���-ɾ�wND�V�Mw�;����mV��U=��ɽ#�n��ARj5ǲz�����@��;���l��I��M��M���'@�K(��ef Y�
���Cf_�dI�?Z?[�d� ���
�/�Z�b\�@���﫵Z5~ZLl�J��xUM�ԿL�Q��,v�@���ᘥ��!�оF��~�c>�:�ᮟ�H=�?��B��ʼ*�'� ������Wl���Vx�9�ͪ�Yy�e;��E�+J;���G�\�[�{//���ב����e}�قe�s`�Wc��d�Sﷲ�I{L!'���B���B)����%"�qcvOO�.���	�s%.�F�^gԬ2������N�s��6��^H1�Xry}�fn��;�i4Xq���p�A��D��p@4/e�V$k+>X�����h^���%}Z�&z^��s��i[&b���R��]�JD\�ڻV�M�ʦ���]�ϰ�6�%bg���ч_6zd[�Rk��2��*��A^o�Gbu��ȏ�����b۵Z-��6�(
��IX����H3�1H5����"�1J5Qx+֘�=8�H=���l�#!���RM�DŻ,R��ňm�R��I�mlR�ָ�;�����،lV6�Q����-�ű<փa˱��Fl�ۏ��ED�{rgu�Z���ΛCW�m��ڴշU1<�����~6��g�7��:ޟ��o�{s��M�l�����{�����+w�v[f.s\Ư\c\���nU$F���}ٚ�X�{�e���7{X���+����4���.�Gw�����
��������]y���fҩ����^M�k�sj���ץ�S����%���=�D&��"��t2���w�|
�{<�L��J���U�ۚm�MdR)��d���ч����_P�/�w��)=�����t�-x��|�}�M��l*�=;�ݗHd�KjT���w�m��$21���^#� 䊓�^��.x�|K���	L�쪬vyrc�$aMZ�a�<?�8�W�Yـ����꘤3��$������U���"<_U�m��lq�S��d8�!���ZS!��l`�	�"=����Mg6�:Q�a��ZiQ[�:�E������_��j1�k(��Ko����_�vx��G�r���_9p�J-K�4F�Y������BZ<�5����9�6�@ZU��bV)w�E�@4z%�'�ZN6/́ۏsb�i�p�=+�D�%竰� ��6Z	==�2����i�S���j�c�Z��#���ʩȇ�η�n�������%���<��o�wa�������8��4�qA��v�+�����K�?!�B�/��w����_�g��V�?��KR���A�F�wg�f��Op~��6�9M�m=���/~��v���B~8eb杈�~$E9�ڙy�9��FAH0Ԭ�49�Nf��Y�����cɄYW_�
���쭐�Цù?��>1Y�Lt�坝+R�?huv`��ZQ8���f������N�)	����c��m���u{�F���eݬ����������W���`-�����d�P�`��_�)a�O�����2���ŴL�I�:�wZ�0$�����sU�?#"1B�y��xU��4ij&/��W�:��e$GBډ.�Q��U_���)FF��:7�h^I����L�Kæ@��.���39k6�S�F�I��沦`��-���뺜V����q�2�R�tX4\ ;��L�l
F�R��4��g���?ˍB�� �V�����O�,N�^�@�'I?a�_ǴO��v���C!:�7��@�w��~ᛯ.i 4Z��֌�t7ckK�&
��~L�j� �X�����N��l��T�$�J�j0:8���c�g�U���'��儂ӂ�PJ 2��˵���K���#]����N*��Z�G˼�ZiwJ r�֚�����[��k�54C�y9q��^f��=L[�����nJ�c-N���V֖�ۿ�-����.�����-á����)�4Q��TYZ�H��J�SZ�����`����:4��������:\輴W�x�y���8�g��dw?���T�(DY�Շb���C��DSb5c����Q��e��=�F�Y����bM�Mu"�[b쀓6#��3'��l�&C�*a�㉫�;�8�����g�I^�o8a3��G������*��t\?_�/d�n�[�lZQr>�m�0p����L��WSx:&���e��2�stZS��`�Z��r��P�r�X
;>7]�a�䔚��L6SdtG�oǰ���<F�#��~�	��Qt\��������>�d͠e�H�Q��A41��s84��²�;�S� �<iۀҮ�vVb���l��x!h \H��t�����YW�I�^��g����U�;P
�C9L�����(�>����k�����j?ǣ���gF�3`��4b���Xh��4�g�Ǒ*�V��K{�Џ�ߖ�ZW�R_�>N�����|����kEq����������S���܂��#�0���tcU0V=�I�~�:��$oJ�!Zu�T��=5�A�&T�X{�H\c&5��w��r�|f���3)����\���I�f�2oK�ں�2��h}L$&�JF����p%_�H+��q�(�C7hr�Y���S��̏�t%�w�p��w��	�&����������Wpg�Z���I�E'��x몯7W���5'�B�g�՘N.o?���Ľ��dd�3��$�צ5Y]C��Q�o��gw�t ��N�%���*̫�O�� EC�h���V�^�u�f1s��0���#h���){{fE�6K�$d2	�rڬ��j��9��s�5����Dg�ކMb%�t�I���;N:�9`6� �u�=���g�m���b"X�3��9��{��{�b0ٖ�M���ÿ�]�D�)�K̆����ɑq�*n����r�vQkZq���C< ��nj�Z���x-#Y�]=��<0��QVn��p�X����{[�81H{x���-�ڟ����Y/��Ѭ?-P���|	%b9���	�d��Ct2l���l��y��QO�6�.Gr��{ޅ8��_X��ל�pj_�91��=��@��^%�vu�W��Ց2��mQ
l�ϣ�QJVOA�5�+c4z"Y�4F��[��Q����J6@
Y�Ga&>�8��w����'�q��V��.�UgG��i[«�=�$ܛO�
O�?�I�4
�/�x��ñH�	�5�F�Zف�u�N���!����"�zZn�����O]`�vXD+Qz�WH)V��	� �6X�b.�C����� �`8j`V@��u�ub�P�����vd!O'�jb�)�J���m�F#��BmI
����n��L7� 3�Zg7:5�,��x���?���l�CS�e�^ ���9�*q?A2��C��)Uh�N��k5�x�@�Ȕ��������~t�lƄ�EYo����tK�u���xl�]-����'��}��U1��iC���ۣ\C׬��=�t^�rrπ�&C{�=]	0��^���+����P��M_��Y���]�Mz�k����%��Gܔ�s� �B�o:�5Y	u�#�ؑT<�z"�J��(`
z��/F��;��U�U�>���Ui^VX�n��j-�Ŭכ-�i�F�4��;���W�x����y�%<:�
"���H����Lt�HQ_��cZ�f�t����07:��Jz��V��C�ʦ�>=3x7~��
V���忙]3T�v��8?�P��oN����2�����Zl�<��l;���ײ��x���g�g���x�N��7��U�rHQ�u akj�w�t�x	x�9����8 F������
~JE�
Oz0z��+�_��X�dd mc=�@�7�S���i����7��{���9;
�e�V��z[T'�&+C:��3�Kԣ7����d�3[=���`_֧ 2wz ���U�+��qa��^�B���v�ZM�94N��@\�6����4hx�S�ܺ�*��n��^P3
%�U"���MP�1`�~m�|�w;}�&�e��/��bfU��d�4>��~���㤿M?ih%~\�o��k�|�~�A��[7��?N;�
�R)m���e����w:y��㷛͵9�h�=����~5��H���Y1;�\ɛ�	�!��7 <]k!�P��@yo��+|<�{��S�9Gv,���=���7�/�3��;t����Y�HO��\��RJ�����z��wU����u\��ֱ�k��"��AGǖ����{W�wm���C	�T�Ċ]%��_����"F�iy���H��Ѱ�0%ی�0�	B���'�z��,/��$�����RU{�r�L5��#�͌����8Y��џ��iD��Gm�`գxiz��C�Y���"e�Y������h�|Z\k�����
E������/�y�֭�ָ�vlY�}�=��&��@W��������OOjϾ;Ʈ��������`�o{$����t焈ߧ+׎�������^L���a8I��"#X��?^Q�O�?�HL��u���`�@+��#�طj�c�g�M.��(��`>P�-Y�w[����3T[��lه3��\��Xw�c�q��G���N�V%&��л}��l^�{���ǣ�D��Wj3��sucǠ!�R�g.hϤ�a��a�������5jAkic_�l�b)m���P���}9$��򾼿-�T����S�u�W-��޺n��^GhxKq�
�����4�q�i�~�Ů�i�h��c�(���9�F�����R?,7����
����Cm�5j^���2�Bq���b9�,0Wa1,x�&7_�U7x���/�ԅ�4�o~��i�L��.�Qsw�wx�nG:dWpr5�I�ܹɬ�m-�û�������3:ԙ4ƻ8��J9�i����]��V���H�������^~�j���b�9��Eq �H�r�`�M�rC^¤�.l���hF���nO)�(��lmE�Ċ�����VU����]�|�Pϛ�toݾ�g�|l,gW3�������͕*�Q��u6�7����)�:N�vy�4Ӑ?c�i�'��6,�l�O6L���u�B��si+�k�bi�7N�,VC�M5M)��pC�)����	��S�R)�dlf��VCp�
��vD�b�=��z,�ŏ�,���H_�Nq�����%��!K!����tKI�iJ���.w�����`���On��ͯ.9�ZA�L.���P��,�<��H�������,v������}��g��yf\܌-rq�K�݃�9�Pٻ!ѧPQ
%�s�9��1��wL$�J��q;����Y7�>��˗X�o�|�U�\�pp���B�뒼ӑIw[��uyAg�8a'����c�	�S?+��k��b��W�z9)E����
��=Y�K��;�+Z�ѠЦ7r�n��| �̘�wY�4y���6��B�XL�JM��g�l�"��Ŗ+p��ko^5�9+ώY�s�W��*�tw�\�Y>\įX�y��J������J`5�j�d��%W����=^g%�.����xs��ǭ����d�ި۫U����1�5Nf��}7\�p�J���1gn<a�5��I��4�=�>gآq�Y7]K��`厫�

�c�P��gudG�c��!?�/$V���P�
��;vn��}8"�;�π���Ѐ0d�Y$A�V����2�vӶ̝�l�,�r~�a�nK���1��\�q�*�ć�|�ж7����Om6�}��nJf��OS���_p�(m:�Tn�{�;�i꿶�3����^� YK9\/���>�L���X�^�<�P䟠�ZʩE��T���CEm���쥊&w�򌶣��)�?�_�)���¬˧���������
��-^{�r=,��^/�PK�/�_\�҆6�q��D��<R��bE���	|Se����M��TA��
(EJ���[�t�ntaUi��m$MB�Җ5�e����U��(�/�:,\�mǥ��(�ŵ*C���<�&i)μ���|��Có?�|�sνwB�ߞ?'$��.X<�1�1�I�9UF��k�G.t�.�ll��rQ� ��6N1���#��erɎ	"���ɒ����$[N�m�ی�)ʔ�)�Sy*!��;�p��q`���b��Iڢ��obr�I>����2m����+��e�3����_�%Õ�,�}��Y����*�z%{�i��nӷ9�r�������{?�������\�r��iO�,����#��F$"��M��*��񐗋_.QC�������+s�渃�\i,��R������F��Wy]�Gι��ys���r�;�s翈���.*X��ʷ������\}�����XYU��9�|�jM�;���Ra9d�����2�[�WV?S�������U�žľ���5EK�]��ֺ���]\fw�{��c�1���ޥ���,�t��ĥS�Δ$wi�ҝK�,��]���n�}Z�j�F�y��o��^hlh<��l�~y��WԮX�b��kWlYq�Vܿb׊�+������Oe��Uw��o��zW�W�2lu��q��W��޽z��5�,�HD"��D���<��?ȿֿv�a����iV4o�V����޲�e�i�HD"��D$"�ђ��D$"�HD"��!i[wh���w��xCƆ7t�f���'��ƴ�[6q�r6�ج�<c�[TT.�2+"�HD"��D$"�HD"���)�HD��
��������؂��E����Z�e0F�K*�X�RY6&��S�U*�����2�ORY�]�Z*k9Q�,�u���x=7W}�T6p��{�rt�J#����鿢�k�&He�S3Je���Ke���� ��ac�8C�v��
kWs�����RY���}*�u|Ip�����T6p��T�V�O��1�E#p<��S��ʌ3+3ά�8��2l��ʪ�vƙ�gVf�Y�qfeƙ�gV���/�ʌ�NN�R9#�¥�T��9��\�?՜mY(y87�4�Ŏ��KBO&瀈\)�j�Z�yi͆�m��V����P�B��k��b�f��\-�\Vnº�tGJ5T?.�i�\y1����D~�;XK���f���X���Y��-���F�����y�����Nmp�V�j�A�f�^��j�����qI��t�z�Z��2���Жz��Rj"�ki[!��;��\���6:���aOB�J?EI#y�H۽�L��E>����-���,j��Zb�a�Of0�=f��(��+�U�G�jB�%=/�B�Au�P�^;>k$RlU����Y��N����S>=�j����t]�tvjc�^�Ūf�_ɉ��vy�:��|ܒ�N���]ٚ^J*���Mma�!�e�;��O��<�hU��f��5'=kٯ3�;G�d�����#C�[D�5�y��%�'��?�qt�:�B�P/Ei8o����'�ٹx�7�>j�gM<����X#��\Z�+�	-�������>və�M�t���.5��Hϩ�j�)Vϕ<G���X%�����{Z�'�]�� ����ɯ����sى;1�F}�'��"�?&�@�@�l��/r��+\T3��i\2�Jْ�u�xO��s�(7Q��^DΦ	�f��˫�5T�A5Ֆ�9��@>�~3
�<r��,�4QҌ�/x��h9/X��M�<�2 �ܒW��i7���[�&��RN�ьb�2��)�?1�4���甖��g�	�]�J�����O�obp���,�@9Yh<ĬA��N#�Ac�E����vgI���}<x�ՙ�*���`wwQ�?���Y��'�[�+��kz�K�-�iAΕ������{�4��Ok)�=s�b��%}2�X����OVz�K���CF:h�?���,�N&��!����Z���g�գi��I6�O2�^�HO�L�VN~����GBB��`�y��>Q���S5�����/YZsq��9^��P�=������Y����(��G����s���=�8��HȻ�t�����w9rr%���=���f^`��b�)�{"��#�}��
�\T#����̯�����E����N�S�\�.�?��
g$d��nv)�[�X�H��N�k�=�N�ƽ�7%O�(�����Ǉ1���!���Y�ǅ�j��g��~�Mf�������-�zEM�N$�a"'����0�n�7}�rP���2���.6�NU<��\��0Y:q/�GP9�����S��3+��4}}:D��r���Q��ӷKF����~�=C\��Kؽ�w�|�2��Z ������il-�����.�~&�'�)}gyi�`gU%�=�=�|����R/u��Y�����z�|��L����Am�%m"�h)z梖��l��È2�=�y�>��q���(�g�h���DZ'�+0�k��&n>�Ä����R�v!Z�IGfd��uRΥY��W�Y�"_�'2M��.-�U>�Q֬�R��'�fb�|�џ�C�EA=s$M3)#�2Y3�i���%WF�Ϥ63m��9�g���d�$�V6��+��3"�@BVeRyT��,�]�����-�w�b�̦��Qz&�����BV��ʢ���A6ʅ���+��L�Ұ����G�C��}��g%WLk�4�h����M�β����y�MtT&��,�!9�{���w�=��4a����E�j�1�V��+��>���I��ʂ;�ne��N1՘�.�-��U��\��c��]�$1��K�5�>�Xj��<�l֤�<[��� �m��&�M,07��}��Uc�����Cf�de�$�b�WZ�Xjv�k�<���,A�lW�S̫�z�>�v��_���g٫v��!J;b���^W��b��f�M�wZm�Wk�������ڦ�^�M��U٬V�Ut�V�j�Z<v71��a���v�7)��Wy�d�X�����b��Z�6��Mb��W+z�|��qa_��Ja��V��N+ x�6�7I����6���c������ś(z���j1�Q&S��>�K:��l���|t����pD[��p��Z��un��'ڝ����f����U-V�k��l#��ч��%�$Q2s�W�3;�DK=���M�9�c�-������z7�+֠�k_��>ZFL2�8�:�qK���l��R[M���	��4y�i���"rS�R'�A�󘭶:�g	��i�3k@�M�-.��ۼI���w<NQ���\�Z��흖�luY�Iu��$LH�5�]5���)�\?#C1�Qo1{�]N Ǩ�f�z��a�㐾$q��Ě�z���8+i& ,8Z�-Q�ڽn80;P�ǎ^����h���}>,W�D�����7.�\�&;$�j;��Zo�%w\���d��Χ��n�Ӭ�ڝG=|?���	OI��ga6+�I[E�u����[�C�P?�ךN	$رb�������p��}�*x���B�ύ,`�3ɘZ��ݗ(�|�'b�qRk���H~�.���.-De	u�Xe�BW�3�)�CH�|��Lj�/��mV�9��I&�d�\,��8^�4�2'�����҈2���l"hK$6��o�$(�$���r8^<�l��k�X�A�#!�@��̈́1X�D1]tU!�9	3MԲ���D!������?gHYN���S�dȊ}�ˤL��x���fCv��y�4��[��nD{��a�����Zv��4����$�۫��6
�]���4`�tU=	^/i��&�p���h���2�iUe�-Y�H�����3�H ��26��ՅJu��f���c8��Nosq��e�����#!Ò�]
c�)R�����l}"�f��l�����8����L H��Ĳ��y��&1�L,)-���m��e��>.Q��_�W\Q.bDifQ��8G�,Z ^�_��(�旔�����R1��� ߄���������\q�㾞�HĢ��"�PZ*�TF+4�f塚9+� �|A���_^D�����bIfiy~VEAf�XRQZR\f���X�(�(���
ME���M4�EE,��,(�[eV@�R�_Vqɂ��ܼr1�� ۄ�Y&h�9��Ķ�QY����bvfaf���*�*�t��ݼ<m�~���U�_\D��*.*/E5V�����/3%����eHNi1�'81��.�yE&�
A-�9!��2SH�lSf�*#��'EG��|-��F�����џ�W��_�Ӌ|=�z ��@����<�A߯d:��	"_D�&���k�&�]����s]
�_�s|~D�/��t)��cyg;>:��j�v��Ad���l��ƒ�Q���s�!�U�v����~��o((�x%~f��s�9�΍@"���LS["&�[��DR�F*5q�HX��h�;��rOpWs�������>���q'�X^����1|�ė����|_���*��/�]�j����/�o�W�;���C����|�G�v�]�1�s>����O�A��p��b�0[�**.*�<E�0_�XX��	�u��J�V�f��&ᘢ]���a�+�SB��p\���C��߅o?�	��<�G%�(�����&�B>���V�|v��s�s|�>����� ^>C�'|&�O:��O����	>��g3��>���(�<����&�| >_��|@���)��g������	>��s����>��g5�\>w��o�g���e�y|>�o�o^�V���'|R�gx���Z�g�\>��'|���*�Y>M�|�����)�9>��W����Q��'	|.�|�>V��O3�� >��g�<>��χ�s|~�7+4��0�M1��]��?��|���|j��>ׂ���s�<>������"��>�����+�����W�x�[H�&�k�|����U�|n��ೳ/ݘ0>�O���O�T�y���O3�� >�����:�|>'��y=g凃�x�>E�s5�\>��g=��>���c��>o�����-�L��W)����>��O>�T��|\�|����g'�<>/��[��>�|>���'a��*��Q09&��O.������Z�|v��.�y|�ϟ�磾|bTa|. �	�3|� �E�|n ��|��3n"i.��O����|��r�� >���>�y|:��M��|���
%�P�]�q|�"|
�g!�ԀO�l ���|v����%�� |���	a��
��B�0A�'L���"!OX-��4�O3��>w�������:��|��U*���
?(G=�$�G�4��~�unA���3|�O-��W�[�g������k�
d�y|"�\>W��
��>w��S�s|�����'>1S���P1��
�aW��|��O+�l����i�9>�ϗ��#�����0~���w
&��P���|���n�y|��}h=>]��� ����ߕ
_)S�ne�p\Y)|�\*|�l����^�y|������gr�ר�'66!!{es�&�רܭ~\�n���h�[[p�vk�������ߧ��ҳ��;Z��iN�Y��(��E�DI�n����::��u�mt����޻u�-���B�F�Nwkk+�H��Q�.5�jkm��T��3�ضJM�Q�����9��Elgg�Θ��_ū�ݚ��V��
���TJ^�&
�i��� :�����7j��Fi��� �T�mm�~7 ��v$S���V'�j��4
Pe����@{{[D*��=��F\tK���;.��J�tPRa
j4*�W)��*�B����]j%�V2e�t2z[�*�SE������J˩���V2�h�COI�&4,#�lՅ��+Lg���+6�2#��/`���U��<(�y\�ҡS`*��WF����~A�������S�Q�l��z��&V�V��4�h,)i뉍e.@�L�IϠg�*=��Xb���;��4c��T�@F�R�y��.V�����x�����/���/Z^������B��o� :���͸�j08H�hB=3�_7�3č6�ת�ၣb�C;4��!�mݤC�i9����ibG����"v����6��ߊ������z���:C��B� |µ��Ԣʶ� -��+0Y ���BH�B�
!TB!D{�b)�P	�*�"n!�!��;�#�P����ʈ8�2��]R	��rZ��!�2�5���㵚��q�f�����xnsK��?��P�G��%�kn��I'�G_/!�Tr�G�㵆 �;2n���������q�ƍ��]Kk3f�%WA�D+�X�%}x�X�Yx����a��T[r_���jN�>+]Z=��&��I
�?	6u�&G��өx��=���t��t��v)�J�tm�U���$O��+uJN���T�W�s�c@c�5�!�$E�� �jCa���E�:��$��Zu<�1����ڰ�;L������T�Vj��$�G���B���R �I�$����.�<�dK�t=�&�H�!��:N����θ�O���u����U6�K��%1٭�:9ق��ĈQ$p7P(Ix�y^�IX�<�@Y� 	�-�(1,4E�B
�B�R��Tm�$��֤�{�>���P�y�J�����zB��c 1��VA��(�#O(�*��~�`�S�z%T%���®�R�2�K��t�P��A�R���:��Lfm�LR՝h�A�����rx��@��J�����׮��y�tv?�"K���:=��T*���oo@�lI��UHв�Ed��3%e�+�IU#��"X�p��Щa"�n���x$�Ss:M0�c�^1-�|�d��ʕ�V��ד��d�ɴO9p(��y ����F�jO~<����?f}��D�h��>�����F���p��
��5��������>,�I ӦPDK!��!M�Jz=!`�:�j�W�����j#(I�8.״�:���ȐN�U���ܷ�%��(��[-p���j2�[.���qz���D.�d����]�?C����Qf� �<��u=�Y�7�G�\��P�~��Z^���*�΁������s�+�s�a���ɪ��]�y��@\ �=�=�-�-�d�u�u�f]5�o��AZ�-�f�Z����'�3Q���0�>h��`Нf�Hd��`���͍-�˨!ǥWs���K�m�n�X&	D��،��e��eP�-b�ز��>/�W�kZ�͙&�F���(gz(?d���r0A4��xs3K�A�^]x�oЄ%���Oů�󚘽�N�%L�{��I��}���
Z���a�eDJ~�Q��ZdZ$^UFF3-���6 ��i�|vBZ��Z�A����H����a1��1�
C�ِ��ܭ����C�+���/sh� �7��!��D�FKr꠹à&����$��k�%m�����@R���#(p9��!C�fg��B[������:� ��O*�r	��>B���Q� �D���
fV&YĠ��.���J�?�_X�5�W��AϹ��\ L*��!���\^oa�>��$G�$����'C'�8:=���`k��W܁x?����A���y�i�ښ��ICo���5�{�k�GG޿���C������89�<����!:�[*��2�4 �5�q������Yc8�h?��)�\'�A��#eV��HfT]�#bT�Íg��ƅ.� �p�>�>U�z�˖��Շ��<Fc�1�H_�Vv�T�;;_Y��uD�w?� קﲗ�j�h��/��^C�k���#l�ى����Ǫ��쩔.�_Ӊke`5f��EGG���VȮ��썎29�����|���v>��}���Nibإ5��A�v}f��#�%.�{��������O�%~@���V��|�Kނ��5�'�[�Å*dn:][�pȋ.�_n,���m�'���l�n��kFw\e\%�������q3��;ύ�9��	C\�nr"Z��sep����T*C:؁c��+��a���6���qrWA�Ѭ;�����X��4�FZ�.����&ui��ՠKo<"�`/mX�	�P	Z�T3Th�\I�<����s�\\�ׯ��ѫ	��h�0�Z�ڱW K��ԩ�*&��e��D�<�D�wQ{��bT]İ@�\��]�_����(�g�TN��\R�����LO�3Q�j�8�\�k	����cC���E�X`�9�h�O������{Si���7�����[�C4�V�7�lA�/��ZUԄA1<�3�U�	*^�7�)xe{�q�11�e�ݣ�#�T��r��G�]�L"��S�GX��[忟�s�s�L�~˜�cW�7�U���f��vA�+�'A��F�T�~��C�4F�壠WUS�P�+*�R�!�`�<�����)��Ҩ�.�Y�\Nk�(�Ң|ހ��r�1����B���:��2���-�deG�N�j�Ԙ��6%}ʤ����U�k��*�E��_?XYX\R�2�x��rf���W���L���hZΔ�����&�g�MM��8�Y4b@���/������(Nh�qh�)�y�{X?�^jM2���ګT-	���}�����;�y\��}oD�>���x��u�x|�ě��`L��s�|�����G᡻����|�f�bXv���r�'��=�!0��b��n��E��I�O����UFw����uv嶥}��z�mZ�_c�zZ�\=6+�������wjh���A+o�~�o��������U��}�ᅻ�[���?���u>;���!�MW�&m�v���]κ���g����w-_�������q?-�����/c��/1��*`��/����y���
qtO3��(�H ����sߧ�jM���[��|.�E�AZ�C#�(�C�C�L��si�[w,��e?�cʞA�r2 ^Yh�ߞ�nZ�%���������%vҚ,�
�79x���!�+�0�8_�A`FE�UY`�m̓�F���m`�ae�q0��"�����4�R ^�m��W��m���Қ�c�������&nL|`��T�5�O\9L��X�z���u�_��r�懢��=�;�lE]�%����_/�m��ʊ�_��P��G�SK�F��v$�ϳn3]p�˻'Tܼ���}�8���.״���S��/�'�w�>�7㴓3�^�+oĦ�MYw_���C�:��x���mh�'��,���2�,>'�|k��w��I��ܻ&7oNN�L�=^3��f�_>H���I�|�1��g��ֺ��9o��pk�_t�R<��W��`m��տ����GK��dlV�HcKc����g�ڒ���4�?��il���,�������2{�@,�����Ҍ�))�F�d��BU��W�O�N��O�Q�'�v�����tމ�+OxZ���[[o�y�C�7&O��4�ƟV�o�[~h�3�K9_�p�?+G~�N�;ڹ���^�IB�wʭ���=uޖc�o��~���5���&�1߳�o3Z��ޛ�6�q��[h։�F=0����|��^��/�n<����l��{�����Zv�=����(�y�;//���Q�G�.9�F���;'�������{�S>Y���w�t�G�{��A�����a��~i�H��?��|�[/�K�y~���=[�ҵ���~��������/�l���,�\D�M��\�ბ*���CoW��Zy��5�_����|�c�6c)�>G�\to����N3٘J�Q�'�N2SR'Xҍ�����'_Z5y���I��'MM�hM��RmNM�2���'�9���D����aii��{�z�ͧO�f(��K� �~/��]L>&�&�i
4���
#�V�R��n g�3l�3��y�W��r�p�<���yϗS|���?����x+p���+;hύzk���=qۢ�����2����������1O\6�1���­�mqX{�k���6�o聧r}7a�����O�(���b_>��sJ�#�^?��k70n���#7�L�'�s^۞����$�̽J���-GZ��>z{�Ń.��t�3o�9/�a�Ɠ�cl�Dsޜ&,LYt�5�<po�[\��?��L�W�}�|x�u��8�u���?xLܩ�}���[�z͝�kwL�S�xr�[�O�:U{�!���X���}V�͊{,o]���~|�����󐍟�f{�����;��.�Lsa��w�t^���V�i����z��۽�ެ%/6����%�_�����������o_z��b�L�'+����3�<���[�޻|��ss�^����<ʵ��fl��e�,�b<3R$d	�}�I��d%f�¡!YF�����o��B*q�-�rP)�;�9r��=�?�ϙ��}ߟ���~����}?���Z��R��yG|N�+U�%��@/�]4��e?������Gc��2_���sGߚ��^������sGh*L���~��Ž�һυ=G|n%�tԜc8z��] ���eۮ�CjI<5I�8�Ŗ>I8A��� �e.	�$,nC b��zhK���a��B�,�˲�#h?;%����}���1V���M���i��CO��9�9��9�)�������a���H��4 Gwr�(���^�w��M�,�L����?R;:֚n �_�t�CW�i���[����;K��8��¥�\�f��SxL�����e��H�����DZ(*syՅ[b��d4�̤�B��QG����lK��T�r?�{���
���QYd�\!Z�gbH?N)�xG�X ��.������z`+{*���H�֤8��WT��~�9�d�ǈ���t��y��Ϡk<�{.Q0��C���-��٥�����������x�7>dT��
h�H����S�Io� `�Qj��tإ�?�.����DEE��H����&���5 6m[��� 6>���w긩(~B�!>1J��Ip�i�7O3���p2'�X���*-��oC�8�������q�N3y'��o�x4u@md�ILL~���d<Lz����fkJ�Ã�w��bt@���V^��§u�T!zYr�NW������������U��_��EU-_-��]�P��k�.��&�Oƻ�k|��L#u�r:I\H������t���35��	��*��u�Vƙ��J�i���Fi9Q;�'�
}��3g�\���� �	K�����^m�9h{�~�&�r��ȗ�r��탰2�����;��ٜ()5��Rd���T��"9�����;���s3��r�~�p���m��~�J��8ro��-?�*�ֳ�,"�c�qg-�UYk��2��l�/a��,6�yJ�Ŗ�=K��Ku��t��f�Do*L[D\S��r�t1(=��O-Vԏf�B }�Q��~��B!���7�_Gc��g3�Y�yؠ=N�sm&O�#XA���J�8�Ľ���A�Խ�������Bb�U���Q0)ԭ=�9Vq��9��/g�=���~���iwk�=S�����jeݧ�E��$���0a�x��	�h���?Q��س��o� l��E�Q ��b?�_3$	�(@Fn���H�\��3�{v��� ��A�¥O��܈�>�;8f�C���g�p�{L[�ߩ���B?m�?0x��KtI�)���]����<��u1唐gi����m�p�QD�����%�t���Zt�⤞v�B��HM��FT���kAP���<�Z9jM`_U�Fֱ��Q&(?ǁI���_�Ɔh^Xc��b�u9���������̼:���`�7,G+Ѷ}��I��W���z�Xg3���L��O��,�6o�T��zN�T(�(M��ؓ&�N�4�_F�Y��1���u����OVRF��[�2��K��i��������
�ɝ<��Byr	�`�m�9{^�8:�.zT��9���a�=3%!ʥ�`+��cgl���k#5E`��@����DkR��4-���R�pb���7����p�zz�b��@x��((L���.�,sm�c�Ͽ�ךD����!.aocO�UHE�2�n]��>���"q���ƑKj1-tڭ�y�R~��ׂ��%`6�R�)�IG��E���]�ZV������et�;�I������y����`*�
�������wPޝ��J#U�R���!�c��p#�����hE��Ѡ�oI^Kr֝����C��0g�s��>��s*?���q~? �M�y>*,�� ؤ������ҟ��إ�.�"��Ez27/{_�ÙsW?/���	���(>
m
��kM�֚n�MƐJ��X5�v���D�e92/�1����E zu�Cr��Ր}b��BBq�ٷ�+�s���C�^�����z�<��SDb�eu}�>��=�Z�+�T.v�mz�)�"�2�*p����	L��v|��,��O��_}"Vo�e��y��>c���+"5G\I����K��m�vu<|��ʊ�����Z�EoᒉR������t8>M�Q��'�%o3�ct�U�U�]����Qq�D���h�沨����嫢kCG���*,b\�}
*���S����8%��3����n�J(�[ȉ�����N7�mOG6�8�G���-��������Z�qP����HH�MS���Zgoo�G\Tu��m���!'�9�{���>���Z�|��&szo�XkyF�҉�2�zrs���>i���k���Z������q��I�ph}yIt�[�i��,4l�M�t���N��rHR��4�ի3 �E�/*Cʕ�ou޴i$Dg��5��<Ѡ�8#�
�鱉�n���rlx���+GUਊ� �M���������#9����a�t�H��3/���Z�"�ݭl��׎TH��m��$,���2,V�q�sp�Յi
爇������_ ��	�W�6��]��6S�@F	����|,Ei���R�DZ%$#OpI���u��CLG��9���&�M�]cw�(!�#Ę��!�nQ������b��]�����v'������Q�l�T>h���l��蟬�t��#���f�>����/�9�fyQ#joP�3�_G��N�E�ai��L�>�� �v�e��]�`���������V\�z�w6ok2�ʛT�7�����'P#��mr�'�8c�R�~żW����1��:jLE\o2���iIX��p`8)<��� q`6R��-�L���ϴ�I�c�IB���H�i�F2mFʠ���w�:!��o��c��mp�ɸ��&e"�
R
�1��8��������k�Y�[^�P��!8�ra����+�.rc�Z�m�d�a['�ۯ�J/�{�(�����HGP�Z>y6T��2�wL�D����.|���Ϛ`.��\ğ���8Y��y��*ڝ3{쇔4*7��'6q�',�=��3����M��]�ڃ7-���OoVA���F�U�xMl+��C�5eP�,,S���N���/n���C`�}*��կ��#fU�iF��ZhW��K�Ė��b�r�ūQ��4��
endstream
endobj
140 0 obj
[ 0[ 507]  3[ 226 579]  18[ 533]  24[ 615]  28[ 488]  38[ 459 631]  44[ 623]  47[ 252]  62[ 420]  68[ 855 646]  75[ 662]  87[ 517]  89[ 673 543]  94[ 459]  100[ 487]  116[ 890]  258[ 479]  271[ 525 423]  282[ 525]  286[ 498]  296[ 305]  336[ 471]  346[ 525]  349[ 230]  361[ 239]  364[ 455]  367[ 230]  373[ 799 525]  381[ 527]  393[ 525]  395[ 525 349]  400[ 391]  410[ 335]  437[ 525]  448[ 452 715]  454[ 433 453]  460[ 395]  845[ 463]  853[ 250]  855[ 268 252]  859[ 250]  894[ 303 303]  1004[ 507 507 507 507 507 507 507 507 507 507] ] 
endobj
141 0 obj
[ 226 0 0 0 0 0 0 0 303 303 0 0 250 0 252 0 507 507 507 507 507 507 507 507 507 507 268 0 0 0 0 463 0 579 0 533 615 488 459 631 623 252 0 0 420 855 646 662 517 673 543 459 487 0 0 890 0 0 0 0 0 0 0 0 0 479 525 423 525 498 305 471 525 230 239 455 230 799 525 527 525 525 349 391 335 525 452 715 433 453 395] 
endobj
142 0 obj
[ 278] 
endobj
143 0 obj
<</Filter/FlateDecode/Length 18204/Length1 58484>>
stream
x��}xTյ����3s�}f�{&�3�d�L Oȳ�ɓG���Bx	�(�b�":���zE�U�^��!�^h�֪�Zmm+�X�m������k������_�~����ά���k���k��τ  `ń����y�	3�k +���{m�����C J> �ݗm��8x�6�� ݥ�ׯX[�p������X�u�ޕ�`��jW�t-�cS���֟���GQR������k7mYqD��� U�׬��z`Ǟ/ 6aޛ��k����?�|:��k{6uq
] �w��]ڵ��Pղ� �|0�q���M�؉r���س~O� �u��l�z�����Yb�����������ן��O�Y!�8�M�R}��l�������B�1I,���=I+�H�@H�~p܍�@���g�r�˩C�I�S�	�9[.�F��2�Nƶ�업WG�"}�W�D"\4�p��u�!Ѳ1T���/ �g������]�Po�?����z�1����?q�C��8�!q����пz/��9c�C��%�����f��8�!q�C��8�!q�C��8�!q�C�y�������8�Or߿zq�C���_�0�g�ǿ��߷���}]��ͷ׋C��8�!��CW�W�o�r�.�a=�S@�2�f�<X�A�"���o���͒Ȼ�<�_�|�{��΅�k.��_�'��߻�@���:��L>K�|M>�܂om���������7�nܰ~ݥk�\�z���{�v�-l]�2gv�R]��ʊ�Ғ)�E��y�'��s&N����fzdwF�˙������0�a�lV��d4�z��s�@n���SV}�*��N�>��]X�uNA�*cQ��:�ܩ���k*���M%���iI���I�r�WV��{�0i�ۆ���ހ�k�,��C�-�{<XAnHYY/��SnP/[j����L�:o]�qR.�MȚ�S����Hr���P�GA���4o}���g#P�솮ej�ܶ�z�������n�R���ͯ�@�֍��S�Z7�*6�Y��=�%,��N�y�wYע6��
�>�~�^M��d��,6�k�q��ɅRV�,
��綝+��4�6�.�n�5b׷������hS�v�Rf3a��ί���J:W˪�[�]Z݉K�Ra�VOZ��?r��PK�ףV;���zW_��mHU���%�r�${԰}V[�1[�ez�d��3�iޘe	�w:�*w�8�6/Ω�%=��.E5� �Z�2\�U���3$��rV_�%��+�x��t~IW�D�-���d��P>ʫ~����\D_�k�c���S&�^�^�zIF��f�mW�<����9��R̨��mѼK�����*�d�C���L��U���'j[>Q}c��4�ae�J��7➨�i��in{���ٶ��\T^:&�q긺6�Icur��rј2˴�U>?:ͩ���"z�VB�FU�MF�����f�4r�Zl�j���|�y��gq8`�G�Z�C!�y2t�h�3b=Z�<r�
pgf�'9T�0�T4YS@��Ų�):c| �y��Ft�P�Wnu���R�,yC��O�OB�:G'�٩6�@[�$�r�L
-�.�Q�}DcJ�n�s������x�zp.}�`��t�!G���Kn�ۧ�緷��t�����Z�Y��BY�~�
���RV�22�@A��SQ�w�W ����
�|w��V&����h��ȧu����eT��21Z�jO�i�(��d��M�>̴�)��\�P�h5E���~,B�
U��8���yZq��*�~��y1� j���X����������3X��6Pؾ��F-iq��!-01?_�o3�P�|�@&4�:��eVQ%^u�w���Nm�n�`�W�1Z�RLsB!/Z���-�2�uaK5�tT��B�8�5cUͯ\,���v�ho�7ƄF�S���7�J.f��ц�7����vZjG�����80ku�p$����p��;�r��d�0Lzg���~���fz��C<t��by�e��e��9��T"�(��Dk<$U��H,ݾ!u��ٕc�F�xGɞ8m�z��NuM�?����½]�6x�Vy�N<v����."�73��X0䶥Q��:�nN�]X�Y9֓z���&1&Q���l�;r'�2��U���O�.7���i����+4�[6���x����˂���=j}6FG��Tp�B^�!bv#*c�>U��~���]=�f��]�z�W�f֚���	�
��l��Í��%�!vo����%�!GH.��؟��n�ĸ&Kr��-u�sh�,�����l�����O]����g�-�>��QeQkU�D�ͣ*z���J�KQ�&O�k�.3��=ͫ�W9Ym�E-�c#Z��]�h5,	� ��}����s#�"��4�b'vR_�����	����\T"��ץ��܄_���3�D8�H����t�~n<��_�Vw��Xh������T�t�S�yX�e`���6� �S��!��L*#�C܍x�I�t��/����\*�M�)ظd8�A�p���k2�A\�x;�nD���J�!nC<�xZ�(\r�]E8����52�zM���fuhف��(�57J�gD�ʣj���ɵQ:>7JمAF���C5I\N2	�SB��pÃ\"�����J�1��+�}��p�#�6��H��^Xc�z
��ᨄX텻kf�w�)ă�}���۰��`6Ǵq7�Aģ��u�>��y��6�;�C�F\��� �)D=���-��i)�)�-��N�7���ȽI�ġ��_RV�_c�y1Ɲc��1ƑT����|"z�W=� �	UP�e�g����W�r�����`M>}TD�6���Ȉ͈���uȽ���D��AD�S	Q�/"���:�#*�͈"=֏݄��~_��&��B�h�#���L���K���9��/���3�PcB9`	��4���@����Ӄh;7�y�Ոs� ގ��if�2�9 /�����F����v+�:t@�%��� ��ny��*���b�%���B�%��oA�%�+�E�%�5�!�߲�ȱ�׾9��� �I�>���9���F/G+]�V��t9��r���<���sr�b�)��9� �m�!�y$��!�kH�Z�$��$�'A	f��B�H)�"H���eJ
	�H�O�`/	�H0��HP&%J�z�gi�A#5l�!�NF��E=���	1=��r
*əQ��F3r������p�<���ex�#�@ϡ=��<��0�F\�x�bQ�ڙ8�۵Ԇib5��m��u�pN!RX�S��ؠ�b���������C=J����t�v�e�9�ZII��尋�0�����٧0��m�v��1z{���ɮ~�wM"�2x�<R>���z��p����>����Պ�l��\���Z�ܟ�N�?t�)���ߐ�<�w�K��~�u���yaK��	�!YS��*u?�z-
��w_��>�ծi�K\��'*X܋9���kwO���]K�J/���]�Z쮌jMau���q�(������:�f`ɠ{ʂ%a�R���Է������z�ޭO�;�	�C�D�h��(�D^�"�	��	�ϾL�I��x��/Q���Y�#"�����h��ZҤꆦ����|o���O��<Y���V-�7���yj��I�7_��G�m,U�����&V��ɾb��ط��dt��[HI��:��Qe/k����3���B�y|z���i~[���K���� ߤ��*f?�9�P�����@�~����a+����0i��@&F=t�?kz"��Ld1#�w_T/�^#�g0@���m0hz<az}�Y�}YY�N���No�|�΋٨����$�EM�Ť �Q�4�U2\�
I���"i�J�Y����Mc*7i=q䬎+�c91�c9�:��zj�~2P�^ľ���6� v�7_�2�����@��-_���4��W���r_Ţo/b�
o},jhi�[����W(ޮ���������i����oh��5V���V��&���*a}����)Ӵ�@s��>ju��t���趝x��M��Wi>\�I��9�W��`�T��V� 2Ѥ�I5L�[����ʘ(�
�s�썉$,�{k��is�fHiXU��"`Ѧ�������� e��U߻	�I͙ߤV��o�^���lJj�h�����N��rV�qc�����1ů����c� H%�l�� �f4�P�-�/���b�Ί� N���I�h�a�����(n��b���њX�w�$c�����&�Y͜�Em5Vn*�5xw�G:	�$��H�<��ss��mK�&c�[��w����0��i£���  �>�����|���?`��`/<AV�p~BNc��`?�U���p�;�lǒ�`>��MR#��{��GPw!\C�DR"�6�ν����2q2Ͱn%E6�"8�_%p\
�I0��-rW�?�a�Ͻ9&H�n|�D>~�-`|���.�Ӡ`/A��w��q<���|�#���8f�r����x�����:l塈9�Z.耕p�)d��"�"G 	�؂�����0<o�p:��Ӑ
�0�3��C�șkG��bZi"��d���/�1]'��BA���	P p��b�ߓO�5�l��#�`E��ɬ?��I�#sH+�H���� b��,�Uh�]��[�������ԥ���XqE|�}�w�1��Le�K�K^'��:��~����������g��­�8|J���%���*���I�%G�1���-�z�[�m���k�����	77�>i9<��#�F
#7�\�kq�߃pf��(������X񑉇, W�s�����%?$���1�����/)�TG�x�b7*/݈�ֻ���(>����\2��/�S�J.���Q�����i�m>�?�G�΅�Na��Wx\��pZg�//�Й�3o��ȍ#;G�G#oC"�!�A�W����g5��N����UbFۥ�RE.B�,!���-y=��<���I�Z�r
�l�.m̓�ZK�೘��x��������3q6.���q\������T�e�w�;�'�W�Dx#��3y���K��������"�%�=�Q�Vw�.��3^����������}���N����i�ѹ?�#'�k��i����V�
��X�͢�t/��^Mi��EWA+�l8��������Z��"Md>����t	�cH*��`���
��Eg&��S:3��o���r���{	��=�~�I2��r����UBx���In��� �/�[Џg��0.��B�����E%ܻp\Bø�o�{�2~�E�*x�]1Q�T��K$?���G��?d+�dNH��Iw���5l������G�>���O��J�W��!r-l��_���V��O`t��+�=H�aTY�1m��!�5�,,IAϹ�bF���مq�GZ�{|!F�W`P�BðB��: �K#�=��Y�F�IvD����{p;�%�G����v�k��	�����DC��t>�y�����I
��'1S%��̇��-�_�wO�{/,���I��G��t��̦}�Fn=��8̍<q#����9�<��K��5V�/p�WB������B;܎V`3Ɵ���u��p���o�}����A����~���AJN��az�2�$F=�@��NR�t2��ɐ�>�<S9[��r֙J�F^�
��|��c��/����J�K��C�_�h���� ;����>��?!L�RLb��h(�+u��<s�������Ҥ>�R�M/q�r����R��*)�	!/��k={v�EG�Q9K�Nb'����z�t��xI�E�J�2(�w�2��w@Juuڑ¼���8�^d�)E��/~�(Y�H�ȁ�>�����bn�^������f�|6��],�#�)����&��_Ag�� �GA/Vm����$Zlņ��WR�X��$ռ��6t?��t��Q���L%&��(+cX�O�~�b&���_���'�i��sEZzG�I�+8����ӧG>��l%�Uo�Y� ��f�P��ԉ��J�]ʰ��\#EF�f�@+$G��36��O��B�ݚ�ĭX,t�A�$L�6�)ZI8�b6�ui�t�j2��2�*-�(�2dk�$��M��#��F4�����f��|:��fll����E�!��(����l�0��1���ܳn�2�s��U�WT^����Bu&��h1r�Ĥ��qI���%{�ÊI���$�݃W<4{µ���R�+\"IG����j?.@��S�����HL�V���N-�:uJ�o���y�|�x�5�M��������>Rv����Y3�������􋖎=�����
��Z���#��4'��!���n���f�^b�)jC��~�,}�m�� F>QL�X��b�h8�� c�??R&0��`b�f�@�h0YA4P�IǬo���Mh�}L�$��?[��F����y�h	�C��c���e~��~pFw����&�n�NK9-�T�R1���e5k:��Ԫy��?F-ճ�E����Y6:�mZ"�9 V�"�F6q֚�h���� ��*�:ݨ3i�as�8�c�i�++�����W���ML�N���|��4�y�y����g[r�m���e�-��D��2�:�6q�zE�e��w�{�����^�Q��AmVk�@��f�%_���l�B(E��d�X�V��S�#蠎!�w`A� �aR�ـ0�����2�eż�DLC8m+1�.#��1��Πmg��?jٶ^"R���H:���a��;`���S1�bdM9ö�pZ�4���s�';X��b��&�&�w\}x��F
���τo~���,�#_�Ǿ4�ziii�4�f�M�ۮ�:UinG��D>��P{	�D^��)��z�,adKʬ�%��$,�T{�ڸ�6t�� ��zYLx��TԦ��"��X��<��x�^;��w������)x���>5�&}��;�7���F��/��'��1���8���Ȥ۴8�q���1���^.�u�IsW-�ki�-��?��(ce��;��b��2��Y>}|���E���}Q9�K1���d��3]3���E�����-֭���m�X~h�>��o�p��v[��n�����Ӓ�:�]����!)9-5#��"�Ή�xz�����LvZ@J��f3�;.2�9.2F���[3|��u��Zэ�w��0�M\�c&�u�Y볂Y\Vf
՜y�5e��H1�-�3#�[όh��տ���V썞���Ǭ��ѡ�'Sb�sev�8�0@��\Y����ؓ�vX'���%tk�qޗ,Pt��*FQ��٤r����%٠y�5򖒖Zf�L-s ZW�����FL,�N��oHMs��iMj*:1���ؑSmgc*�<II�	:=�>���d�G�׎�����졡�/_�⫳&,�(��O\�p���m�g����<4�/�ya����gg��<��\K�If3WT�u����#p����N�i�~���lK���"LI��ZH[���V�eB��;��u�����q�K}o�{	�����^�	wĝ�v��*�*Ӛ�ֻ�p�'�,��r:��D,�	3\�����t�'}A>�J$���$8]&���.Δ�A�3�0�B'KA^s>��"F�o_�6�ͳ����c~j�S�Zmْt�N$�b��[1������`^fg�;s3��j�T�����eb>f�J����}�\�ݾV�&���8�1�vD�{_�#K/��X�`~^�zPT\��n}�~���g�q�S�o�3���a�7kQ&M;)S3���q�~�,��g�qю���u��$��a<��좉q�������\�b\Ù��
F���kLz�v��W9ʴ��g�Λ��M)vL-*LJƛ4IH**Ԝ/SǕ����ͫ_��sg���?7_���+���[�|h7�Bsk���F�x��?��ˇ٭g;^V���N���U�#O�|1_����x��.D�e��`N$&�NOt`4L�C$b�<�������a��}���l�J.M->�~!�18��/l�F�=��-7��$vb��'�l��˄���َi���J��n�'���7�Mu��/�ee�����jgc�F�_��Dg�t�07��N�vzaa�*J���M�3��u���?�ZU}���ڊ�	�oφ�収�Vݹ��kh����%��^ʳ@�)����z�O y�dC�g���q��H���:�����/v]g��[u�;���ƳuĿ�����ԑ��:���u$X����l|ǵ��-�xȃ��i�6���
X��6xA�^����eQۖ�J+�o��۹,��f�^�c/���ܬ��J��U�� I)��3/۸q����k��Zx�jGҼV�+�j�'sq{FZ����W_�-�4Zs&O�e.������9v�]/���cG�#�
�a침鑼(�^��_��5}�@�7��3��1:.F�ctT�� !�P~a>���G��^�/.ο�%�d1n��ቢ��":��g�X�nL�̓�Ņ��2y��F��S�|7㸝��cn䍢���!� ����laޔ3ӑ�^~~1�cJ#zd>`�~]�_<��'��@|Rx�a�R���\^@&���^��%��Hcjk*mH!��r�����Y$�O� 6�l��.�Ǯ�H�t�ݥ��a��EEyE�$�Å�o�������O��L+M��gQbQWT�A�c��������.ܼ��{h��
l�>}�M�����7Ϻ4|��C(oۼ+��f���[��΃+������5��u�uk.�������;WOv|��o�7���\�,5�z���ϒl���lɉ� �"�~ј�0�Î�U�0^@:��9���`���))*��S����ȓ$�xF��`D�x�݋��˾�=�o���ɑwG�z�h��5��Z<1��+��Ha��hWٚ@�Ȍ��pd�\�9��{L�2Ya"�&Ҁo8K��Kt!$��)�M����v���`MdkÓB/�QAQ	aBP���bא��$&A�
�(����,�kG`��ۺ��e]k_���IBP׻�������?��򞷗931R�v�L�f4�.Tj[S�.�nA��9���m�	�bn	�TP�e��4������j�����;���Y?f��=�y���Sۀ��`������ҷRL)m:�S�:���k��x�K[�^L��)0w��E�E��c@ⶠ�������Xg;��Zv�\�\p���e'g�.�%nI�ttpp�13��}��)PXN ���Z#���W�Pt��\�<�Ы�E��S[�;Y�����\�ч�j/�E\��e���C)=K�-�XE	�����}$���_T�Dg�SS�<<ݵm	����Q.~�h+u���_7S�7�Sc36c36c�����i]������fjc36c36c36c36c36c36c�;�|����m��fl���7��lq_�]�t76c36c36c3���a=�1��Rۣo��Я`X��S1[�2L�����	�>� �s���M�Oھ&�Øc�Om��nb�����M��G��_��S0�Jm���94j�4���ym�n c�Y;���M13Gݷ��0��s�_��[`G3m�ƌ���N��]Q���\���)��������?�- ���k���>�C�O���`H�}R�d�Kw)��I�}R�d�����=�[�oy�C}k�y[���Q���C��=��	G}xG$#�w2�o��&�~D���j �f���I}vC}���>ҧ������u�l�p�#0z�X&�	�����ǔh&
�T�߅`^� �`���@�1>���5��$�S�G�w1��-�����3<�]������ w.���
�S��@_�J�������X �uՏ�1�A0(,�
�C�eka��Q�����G�^&�)�C���d ]�X$��8+D�h)#�G��GTr���G wثB3� J�4��y�=��'�)�'G���K��4�����r���Ѽ�@�)�l��k R�S��F��D:)��'�bD򜍤�����s�-�B���!:8��H�^o�X*ҕZ/O0�}�S�����[���������~�l�h�	y V���T+�/ҽ�#E�J���T#�$!OR�)�!xo�ꌅ�b!��_z8�;�DR��f ~5�~��q��H��4z���y�>�I��#8����rDG��&���X$ڱ�V"	r ���]��=?��F����3z�q�o|�%��3�~㑤����\�byHO"9_�Y�VR)�)�]��{�G�z^ ޻��~;���[�H���
����t��5	tԿ䫧�@IHY4��.7�P��#����F�2��/%%}O�«��Wh�I��>�AJm&��ꬩ�!a�����Y[��L3v]�H�ZV��(E1���^��D�f�R��^�@���X�_f��#�ev(g�4	�ȐF6�[dU!����5?-�a�eIom�6g�^c:n��:�7�>���x�U��#�i'��HP͔i�E�w������\�>r�W��I/�hie"_�k��@2��u��=03��I;����+�6��` �\�)B������[�5$D�+�5G�?�h&膌��kU5��g�t<��m1X�ZTt`mo�Q����3_��|(�J�>�׳����绡��|j(���櫭�i�D:2P�W *����C`�"-�ؚ+,�u:�E��T�z[�҆~Z��Q���<�⺥/�}�VxRJ�J�ҧ�5������QW�ՠ\��b�i6�e���7�1���H]���"�F�8_��&��tU�Y?�J֬#Ü�r��
�V�Z��^s�aQ�^z5�R9�NFYy+�����q�*��4P-�h���u+���Q4��3� B�]�D�JCu(���G����D0�r\��1��� ����#�M� �w���-�fR��cQ$�%�]�i����$��`�Kؒ+.���,�� �v�ps>�?����z>c����� f�3
p�Fp6|&8��F2��&"b�:)q )3���pP?��h#�_<h�R���7����I�s�?�&�
�;����=�VgP�x4j���T�j� ��+V�;>z'y�`k��4��E��־G!��Ј�F%#[�U�֖|$��TӐ'rI,�{H�^�{�w�4x����my�y5��!���S���R/P�l�ȗ@O��037��+OΒ�	
�B����Q
�R�j�
9g�d8_���Q�|�Z�%3q�8I�J���y2�/�W�jp�"S*�E
e�
��!z" �
?�8_(Sf�qB�H!��}Yr<.W������j\f�'C��#��2�H(õ��Պ\�H>24yB�ϕ�%*\��&��R�D�����	.�I���1.#gq�D-RI�P@DC,��25���B��ר�bI�P��+2�Z;���N�$3W&T�^	R�JY�N��ԐL0� PB�R\�J�'�g⼌����R9�(e)dB5OjTR�T��HF5�
��S�չJ�L
��P�5L|�"���@N�(��5
\��5.���@�\(�J��� �|
ոR�ʑj4 ]z>ҦNg� T��u2 �D:׳�T)Ĺ"���2� X^�̀�<@T*�r�бt�+�|�K�M�� `�����>U5�4S3�]��'Ҁ�P�Hr�MUR@U�ȓ�BqK�	IU�( )�QWK��&K"S��(y� �ɒ�K�L�X
�L�\@�j�.T^r�;�����({��I��<i�T)K�L�*��� �0��{�"�PC� ��G��"�"B\�j� 2A�HFId ���[�2Te�h��I��Q#�rH��L�hF��3T 2������L 3�1��(؎+�ADʡR�(�����K��
9�?�
Qn���z�h�bl!-.Ц�ވ#���_���,8m�n��A�u�2)�S�6ĥ"*���J��sbi�� �(s�@�,� uz.^5��z	�����0@[k��UVɀ$ɠ�j1�������0rUr��!+@�E����4:k�c��b)
�����$U�?2�d�fO�.���@�tI�������L0��%�[
�������46��sx��ʍ�D�l{2�4nr/%|vb� ����}�����?��p�&$�s9`����M��#��D(>\� i2����D���GŁ!;��M��c�ɉg@�Ɠ��dnTJ<��'��x �&rc��
'����T��I\ǎ�G��)�{>�/��4�ύ�K��x��0���#�9$) TT<������	�X��X�L�]ZMzl�7*��K�bD���`� R��[Ӹg���>���;x	ؗ�!�@U�-,@�8E�i�%�Î�p�!0\�(�	�W��,���Sl��c�G�%ݺ@{��3��VN����h{i�[<	���>�����ﵓ�K����w�o'�g��n��n��n���y67�woy�]��w�w���a��N�BT#t�Ft���8�JZ�a�)�ޑ΢������{(������|�E��T�0�?��V��qh�?�a�<�R��(�O/�mn�L���;��~8xub�r�<*_%c�*I6�j�l�0����̑?� /���Ӂ$纈(r�gjѭ8���ŌZQ�Z�&P)�aaj�cK��7�����)�N)
�R���0�qYձ��%ZR",�����W��;۵q�<r��������KK7V9�"zQD�XA�R�T� ��
���Q��<�>B�蹥� ������=5E��'ZÁ��e�P�%�gjr�a'����q�B.fu$\����c�t�',w���읛ד�9_�F��ē��DǶ6��D(�

	b��!QX��pfMX�u+{���Jt&G��YBx�5Y �9��Q��/ӝ����<._�G@>< �(��K1�hE�V���Q(ز�a��y�VC�|2]�1��Rv�]e3YjW���n��{
�\C�z�,d�Q��AE5��>�2fN�sr��	����yrR���L�S
"��$�ؔ���I��LW��k\�,���?�;�ν��'�f|x�Zɏ����̏1�}���N�w�>�c�p_i�F<n��^F#�ʽU'�^�?����.�\[^��뱥#��e�8�n�;ψ�F��8�E�5NtÉ��nG�(�0#2j>E��vn1_Z�Y���*��e�h������S㬾�݄�;.���)��(@#&�+P��-݉�p�c������-i�SY%�uz�f�A�tg©��#��5~�Ҳ���Q�v�T��hE$C 7zї�V�Vp����D*3Gg'�H��̖�Y?����ތЊȈ�'� ��oj���ČB��}�8ݘ����������5�=�z�%���p�A/�
Lήj�1��~|���m}N�m���vz����/��X>ޮ)(d�������ܹ�[��=����~����*n��y�S�n}�:��?'��h����v�g�!�%jˆO�w_��n��kV樉�Fl�;J���R�}i���3g^{y[��em�Ҳ�aJ4���u��N���ܔ�gTЖ�߱���U���5ֵ��4ip����੥b������0�zA��!����f7�*ڄ�L�ֱ�.J����u��T�Gԋ�g����ۭ��	_p�:��K	QdJI�A��_�zLa��O(��j�
$�	�H��"��A�f�.��i&z��G�P.&BX,�@2�5	�?v����2M���s�ٜ�|��]��WMc�}�z�ҘݫO+����8o��q݊(�Ɯh��v<�a}٫wt�gS,?u�W>���t�������-zt{���&��_B�Ɋ���p,n��9D���Q�^�9坛�o�Q�)xS�AOG�U���~��y/��8�������5}����s�^��s!�]�O�F����G#�OL4��ծ_�ŧXC\�j���l>�[�����S^^.o�6{ݝ�mk._�J9�!n������q���t^�m?(8>I�=��q�����G�Vu٨ hd�n��t�����}���Չ���}�)�����6�_B��rk:�Ekb	ˆ�"+=���g�phb��@,Q�$��������t����!��
��H�qr��$�Eߵ�+g��\ꢿN�_�P
�eA�.�����;����DJ�B��B�k����tY�$4�5dܞB�D��g�L+�R0S'��iG�<x�������é�?}�!�I� �5�Tw�ѭ�e�k�u؄c�ky������{HM���1�����Sl�²�.'-�-w�&6�u:�7v�K��+���Mt���ݩ�Ev��l��0���7=]�d���3?��j�*���ᗔ:Ĵ�qf��h�����1][u+���^����(�Xmwt�]s�~�>Y�BG�nX3-��K�n���'�w%����dm�a�珯=����V�OO[�/�5b�tRe�+9��)�>��Y���c�C�����O>.�ٔ�9�yWܔ��gߜ_��CɽY+�:O���hAb�{����8&�Jλ�燐ٟ�7�����>6�L���9�dSU�=X�n���Cߋ�儛�7�z���{Ǟ)M]3���6������Uǲz�.^���;z.��j��	��<�9Ux}Œ���'��������"r��n�_:��y�Ǟ/���M���iwq�˅ǧ�<+A�}ߡP�� N=�;ߜ�Gfw���]f�=�(0z���y֣���]���Sgǽy|�z��
3P�E�R��r�����P:���ߵd�3���Ή��Վh�b�B��}ȼٹ9o�
�<��J3�"�F��s5Y
�T��;L,�� "$wp�߻��W�}e���������e3�5�u����GҖ�7�;�����s�[4���٥�E�܅"�o]2��������J�Z���/yRr��D@�˟��ta�{o��{��+k<�g�圱8;t�٪H��7�d2�x�#�*>{�+�鹹��·�Cc�1w.!��| ���ˋw��x������wr�;9sW�a}b3Z{zglX|�ia�Uo&�o�`Q�rrS�菔r�$�)�Ӵ���}u��+�u�f�\z���B�.W�����n����7����#��.�oYO��g�>��W�.a�vmE��+&�L-�5��g0�p	�����
l7���n���-��YS)Z#��ݳ�.�Se���[���_��3%DY��CQ�∿]�_V�0����lP�"ڠ ��;��P�(�߼��[<�v0-����;��]?��/�R�Ԍ�cm�����s�0/�Y53'}O�D"n�TvcL�[i���/wit�o�7�ٌ��zR��up��Iì�[O�7x��߹7kĥ���>3��B�?�[�N�w��3��i���r�s���ٖ�E{*C�e����}�>8�i�<�Y{�7'Y}F��|TV�a��X��<b)���ʞ�gL��������"�^��� ��-<�������OK^��!��_�{o�����r�B��������yL���UK�M�ڧ��V���(cߙ�w�<������=��#=�teՋ?s���(��;vT%d6���T��^���=����+:�����sߋ����W��v��<l�����~)[~���@��ƴ���--��L��zDXI�(�Ny���C��>i��0�_����~3=�eX�:����m��=w���:.�9:��"���ya��ћvT�涿6�}n'?���A3��x<����y�������"Q�X�o�6�&�~�i��'��A��&t����oE3�)����D����$]W
l�'����ǀ�i�H*�'2 ��N@6�X�l��A�d�莆,��'�"ꗵ�
k�s���Uٹ0�\�Wd�������WFv�}`�w{LC�ӹ{'�Zw���c��VOB���V5�^�8�"/��䋧NX8��l�
��YC��\*�nɨ�vm���1ۮ�8>�����Q�����<�̎��C��1i������y�cp�Ӌ�����7��A��U�Z�^����_�l.�_���gs��>��°��n��sKH�Z5F�k���C�65E͛tm������W��{	or�g�~����5������v�ª�o�2�������y�A]jC�≂��Zmi�1�ċ���Y��=9�?4s�����5]�9{}��+�˒�>�ό�����c�ƌGB��^��æ��2�{�p~ݮ��δ'����q[9�U���������Eîv�q��Ŕ��B+[����w�=�s��V5�Wս�7Ŕ�?>�v}ҬG	\b���7Z������[5��6]n�{����k����MO=l���+i����zڔS�5�1�w0��qJtI�E|�ŵQ~�E��G���C�/*�L��jZ�_V$�(��S![r����f�kg����R����W�%���t뎖� =?���-��E��ģ��Ae͍���$������s%��@�������������[� X���aD�0T��9>�D$��ȿW澁_C�������D�B�p�^ILQ8��Б�R���1K���d��*_�T3�49Do=*��w��1�3���0���|��Fj�Cg���;w��A,�Y��%�&�g^����Ԫ�u�h~Yd�����sk$Ø��׵�s9�>����x�C�W?�^��v����g�$�\��?�|��.�{E������};܌����k/�r�[z��Xt��1��ǯ���4�ŉ�ԘnG���[���ziS��,梊nݲ�sEnR��%�w&�8<�y��/�{�=�X�e��m�Mgo<��V�xI�m��3��n��η�����b'7��G�#?n�zw�����q�����l?�����_=p��J����5��ML�Q�y�E�'dXޑ�q�D��x��Qw{w����O/�uu_\|�篟9U�{6�Z���CD�ۃ̖M7�3=gZ���pP(����;��d�����ߣ�V.��]��90���}���
��b���K�Fp�:�x~ժ�c�tz��mӻX���+^���w񭇹��?z\������Y��m{�~�C��Ҟ��M���7o��慝[���;T�֩rtk�1�ٖ��6�\3��r�Ҵ���q�Ñǖ�dY��!é����j{�1I�XE�*����J����ۅ����T���ub����ydŲ%W	��tHm�v��٩Ǜ�~���b�f�%�[�Y�DrE�������w������Wv-�������Td��ʬ|���L/�`~6w�:&��T]Y����l�'����=}�n=�7�m�Pr���eZ���z����u?�]R����SG�iZv�m���X����
��g�6��L�(�����p?����⩸��;?;$軴[�7Nozr��35?̟Ӷ�����I�w�2os��Q�_{v��c�®�O"n�=6̇�]��4�����Ig�5yL�r�$�.����.�ܫ����7��>l����!|�
��C*Vl���B=7�F����	�-7��8�M/� ��t����"��<��l#SV�L�F�9��v��s6�B8��U��B
 �_1a�B7�Y�`Vh z��Gf�Oy{`�Ɲ�6�V������ώL�WD~�&�����&��z��o�y������������a���ݴ��ULʉj�Z�n3��g�v������j�J\bܨI�KsG�\x`���&��!&O�&�O�,�-رn����.�;�޽t���z�ĝ���c�޾��P�5�WUE��ܬ��\,~�v�Yi�6��C]^�P�;y��ݥ~���s��u6lׇҶ#W?0�ܳ}�x������+���&��V�8|��d�ɝ�6op�����g
��vI�7y��K��O��<|�,'����� �O�S�
endstream
endobj
144 0 obj
<</Type/Metadata/Subtype/XML/Length 3056>>
stream
<?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?><x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="3.1-701">
<rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
<rdf:Description rdf:about=""  xmlns:pdf="http://ns.adobe.com/pdf/1.3/">
<pdf:Producer>Microsoft® Word 2016</pdf:Producer></rdf:Description>
<rdf:Description rdf:about=""  xmlns:dc="http://purl.org/dc/elements/1.1/">
<dc:creator><rdf:Seq><rdf:li>BiServ</rdf:li></rdf:Seq></dc:creator></rdf:Description>
<rdf:Description rdf:about=""  xmlns:xmp="http://ns.adobe.com/xap/1.0/">
<xmp:CreatorTool>Microsoft® Word 2016</xmp:CreatorTool><xmp:CreateDate>2026-01-07T08:49:12+01:00</xmp:CreateDate><xmp:ModifyDate>2026-01-07T08:49:12+01:00</xmp:ModifyDate></rdf:Description>
<rdf:Description rdf:about=""  xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/">
<xmpMM:DocumentID>uuid:67BE1923-0546-4CB5-8D78-E95FEF8AD87A</xmpMM:DocumentID><xmpMM:InstanceID>uuid:67BE1923-0546-4CB5-8D78-E95FEF8AD87A</xmpMM:InstanceID></rdf:Description>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
</rdf:RDF></x:xmpmeta><?xpacket end="w"?>
endstream
endobj
145 0 obj
<</DisplayDocTitle true>>
endobj
146 0 obj
<</Type/XRef/Size 146/W[ 1 4 2] /Root 1 0 R/Info 20 0 R/ID[<2319BE674605B54C8D78E95FEF8AD87A><2319BE674605B54C8D78E95FEF8AD87A>] /Filter/FlateDecode/Length 328>>
stream
x�5ӷNCA���d��l�@09�ɘh��9��-�����GB�D�D�d��-��H3:ͬR��F5�����
���#����� �-�n�Y0���`��{��I���Π�R*NO��8�38�c�����ܡ�N�8��H�$H�H�4H�0�%�y���<d��`�@dC>�Bؠ 
�EP%� 'x�n(/��ʡ����j�����ڡڠ��=��������!�1� L�8L�4�`
�`fa�aV`	�aVa�`6!��؇]؃#8�]�|�����"x��ބ3�pV��k;h
endstream
endobj
xref
0 147
0000000021 65535 f
0000000017 00000 n
0000000165 00000 n
0000000235 00000 n
0000000508 00000 n
0000003569 00000 n
0000003738 00000 n
0000003978 00000 n
0000004031 00000 n
0000004084 00000 n
0000004216 00000 n
0000004246 00000 n
0000004407 00000 n
0000004481 00000 n
0000004722 00000 n
0000004998 00000 n
0000007825 00000 n
0000007995 00000 n
0000008247 00000 n
0000008523 00000 n
0000009076 00000 n
0000000022 65535 f
0000000023 65535 f
0000000024 65535 f
0000000025 65535 f
0000000026 65535 f
0000000027 65535 f
0000000028 65535 f
0000000029 65535 f
0000000030 65535 f
0000000031 65535 f
0000000032 65535 f
0000000033 65535 f
0000000034 65535 f
0000000035 65535 f
0000000036 65535 f
0000000037 65535 f
0000000038 65535 f
0000000039 65535 f
0000000040 65535 f
0000000041 65535 f
0000000042 65535 f
0000000043 65535 f
0000000045 65535 f
0000011125 00000 n
0000000046 65535 f
0000000047 65535 f
0000000048 65535 f
0000000049 65535 f
0000000050 65535 f
0000000051 65535 f
0000000052 65535 f
0000000053 65535 f
0000000054 65535 f
0000000055 65535 f
0000000056 65535 f
0000000057 65535 f
0000000058 65535 f
0000000059 65535 f
0000000060 65535 f
0000000061 65535 f
0000000062 65535 f
0000000063 65535 f
0000000064 65535 f
0000000065 65535 f
0000000066 65535 f
0000000067 65535 f
0000000068 65535 f
0000000069 65535 f
0000000070 65535 f
0000000071 65535 f
0000000072 65535 f
0000000073 65535 f
0000000074 65535 f
0000000075 65535 f
0000000076 65535 f
0000000077 65535 f
0000000078 65535 f
0000000079 65535 f
0000000080 65535 f
0000000081 65535 f
0000000082 65535 f
0000000083 65535 f
0000000084 65535 f
0000000085 65535 f
0000000086 65535 f
0000000087 65535 f
0000000088 65535 f
0000000089 65535 f
0000000090 65535 f
0000000091 65535 f
0000000092 65535 f
0000000093 65535 f
0000000094 65535 f
0000000095 65535 f
0000000096 65535 f
0000000097 65535 f
0000000098 65535 f
0000000099 65535 f
0000000100 65535 f
0000000101 65535 f
0000000102 65535 f
0000000103 65535 f
0000000104 65535 f
0000000105 65535 f
0000000106 65535 f
0000000107 65535 f
0000000108 65535 f
0000000109 65535 f
0000000110 65535 f
0000000111 65535 f
0000000112 65535 f
0000000113 65535 f
0000000114 65535 f
0000000115 65535 f
0000000116 65535 f
0000000117 65535 f
0000000118 65535 f
0000000119 65535 f
0000000120 65535 f
0000000121 65535 f
0000000122 65535 f
0000000123 65535 f
0000000124 65535 f
0000000125 65535 f
0000000126 65535 f
0000000127 65535 f
0000000128 65535 f
0000000129 65535 f
0000000130 65535 f
0000000131 65535 f
0000000132 65535 f
0000000133 65535 f
0000000134 65535 f
0000000135 65535 f
0000000136 65535 f
0000000137 65535 f
0000000000 65535 f
0000011178 00000 n
0000011610 00000 n
0000074514 00000 n
0000075076 00000 n
0000075404 00000 n
0000075432 00000 n
0000093728 00000 n
0000096868 00000 n
0000096914 00000 n
trailer
<</Size 147/Root 1 0 R/Info 20 0 R/ID[<2319BE674605B54C8D78E95FEF8AD87A><2319BE674605B54C8D78E95FEF8AD87A>] >>
startxref
97445
%%EOF
xref
0 0
trailer
<</Size 147/Root 1 0 R/Info 20 0 R/ID[<2319BE674605B54C8D78E95FEF8AD87A><2319BE674605B54C8D78E95FEF8AD87A>] /Prev 97445/XRefStm 96914>>
startxref
100544
%%EOF