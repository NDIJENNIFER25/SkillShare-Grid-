conectix             0�.pycs   Wi2k    @       @    ?   ���Q�Ĝ?Y����v���                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%PDF-1.7
%����
1 0 obj
<</Type/Catalog/Pages 2 0 R/Lang(fr) /StructTreeRoot 14 0 R/MarkInfo<</Marked true>>/Metadata 223 0 R/ViewerPreferences 224 0 R>>
endobj
2 0 obj
<</Type/Pages/Count 2/Kids[ 3 0 R 11 0 R] >>
endobj
3 0 obj
<</Type/Page/Parent 2 0 R/Resources<</Font<</F1 5 0 R/F2 9 0 R>>/ExtGState<</GS7 7 0 R/GS8 8 0 R>>/ProcSet[/PDF/Text/ImageB/ImageC/ImageI] >>/MediaBox[ 0 0 612 792] /Contents 4 0 R/Group<</Type/Group/S/Transparency/CS/DeviceRGB>>/Tabs/S/StructParents 0>>
endobj
4 0 obj
<</Filter/FlateDecode/Length 2728>>
stream
x��[mo���n��a?���p�|Sq�"�����ھ��hje1�I�u}gf�/�Hk/D%r9�yv�gf����.��w߽������󷬺c��.�v�����������|����Y��*`�<?��O�:?������_9���Cv�9?�p��8K|/B�p�Kbvs��x����dwt�������Z�����F�g�2r�+��?��f7���}�;����}����C۹m۹{��v2Y[�N[�Ƣ`ޛq�z<=��{:��������;m�r�OV������V��80\ʁq�%�EW�/_��y@?��� ��E�򴵑}��^�Yk�ؾE1�2cQѰ��6�tSG2�ˏ������u[S�Es�^�6(�oP��E�����kF�۹���]ٶ2����o�U$2iRx�3�!���}uNS�`��㯐?KJ�����r�qrg�/w�"��d��wX��ߔO�:w
�c8�ox!��E�]pD:����:SI2o��Wg郿����	��+�_��B1E	�܋�;�s� ��:'hY�;�P�[6���/'È�[ �1��
y���3
�0��_VM� �Vx�1ߺ*��W��S�}���-���<�3��6η��^2�{8,�ǁ?��|ߴ(�y��Sv�h �)Q�r��JV�nHJ�q�`�@����Kq��0��=�)�4�1p%� ·ǹ�=�q�8|�ܠq��h�
�O-�"��)�qI'��k���Lp:.֕G_���� ź��H�V�Z�S�S%�Y1H�]p.H��h��J�������-`�7MF�AEKŇPF�����wn�\����Sc�ﻌ ��ir�� )���5�De��9�92��a&�Gq����(��1dX�U2�I�{�R���n)��a��C-r5�KW�'nV@�"�Pl���k<!�1Q�5�MmAQU��r�'�yw�.���
��+���t�~�s(����������r��1b�x�!��>"�W�� 2֥d$�Z���Im]Jv`���,�Pp�Oh�Q����B�����-��"��=�'\��3E<%/I��d�W^PFA����!�e�ʡ� lР+�ەq朸�91��x���ZC7�[�-�j�L�g�DƾX8VGӑ1��RZUt�'����g`�u1�
�ğ���aK���O� 92�#b=��i
�	8tzf�k��"�;g���R9aM��L���*!T:g�ٍ�S�n�opV?t��y�I�&=R�J�J-F�q�f}����T����5��0�Ĕ����j�1��xȫ��{hW��j�QK^`�|R�`]ړ*v:&�%��xQ:�,%y�XL!���!Hը�Y�Zx�ʡ�Rv+J��'� (p�ǩ*VjZ�OD3T6+ڢ{ʆ�Q�v6�H顺ԣD���	?�}I�9�lm����	�3�7 �XJք!���!Ի�hH��	��W�t�F�Ygx�C/���톤��f9Ճ2#}?`�+�'�ʬ$��jڢ�X�
�������^5�z��"���5��'w4S�.�
���2}�2���Y������X�)��{*��1!��ϸ�TtDJŝZ�#�_����s&DKYɶ�:�L&LU&���cU�|r��N7 ��"`�F�i8P�3�挧������U��`�����XE�
S뺤3)��L
L��Kp�|�$/Y'��K��z�"k�Ӂ�2�zs��S�Mq�6�>{���9�M��T}.�h*�����Ȱ��:Jܪ-���{?t�&���/멟�P<o(��X.��>�x���Ԫ"���M�aɠ���
��Lkj�5�!�]'��4?(b,ǠT��@0�+���$3�Tν8��	F��� �8�,���q��_�����V\�륗 ���t� 0�D�Zuj�)�6���:�
���9�$~�yW��^c�R�ē�B���K�����j�Z��Ž���f�u_R�((����,��Z��˳FȚ�ܕ��&G�������_�9cX�ֻ���M&
m����
I55�l�N'��F=��q�.>��sq1��R���L�����G�%Z���LP�MG09m/�+�Ԅ�����
6۞����ܮVX�U���m�~��fօBjk��"�I$�����h�Ⱥ�B�'�.��,�7](�ֲ�qg��x�<��6^G�DS�M_�^����p���Qj�
<�N�1�</M�-0j�a�b����X��Qxa<�XD$|%p#�s�h����K�v,�[5����[k��Wj�,/��u�%��z��'M9j?M�`�(��&��M
��Fo�����a-b�ir�h�����K��6JE�U#�E�ٸ�@ɺ6����ƹr����O�c�t�,�oq�S�=N1x4�/����=�����x<L�  ��x}�o+uN�r�Z�o��X�"#ƙ��GJ�F�<�phU�'�`��-9�������DLr:&YJ�� �VGq��O]�����1Q���Ma����~}ѕ�Z!��-�����6�4Z�pl�?�\��p��ċfbd��K�F�O2�3y�	Z�bp�	���H;����__���	�м��l|�oM�?#R]����[m͍G{�	j��s�M��!��s��1��}��鯽f"c���c�{+�ؤ��P�?���P/���g��EWF�sO;����i�
endstream
endobj
5 0 obj
<</Type/Font/Subtype/TrueType/Name/F1/BaseFont/BCDEEE+Calibri-Bold/Encoding/WinAnsiEncoding/FontDescriptor 6 0 R/FirstChar 32/LastChar 116/Widths 219 0 R>>
endobj
6 0 obj
<</Type/FontDescriptor/FontName/BCDEEE+Calibri-Bold/Flags 32/ItalicAngle 0/Ascent 750/Descent -250/CapHeight 750/AvgWidth 536/MaxWidth 1781/FontWeight 700/XHeight 250/StemV 53/FontBBox[ -519 -250 1263 750] /FontFile2 220 0 R>>
endobj
7 0 obj
<</Type/ExtGState/BM/Normal/ca 1>>
endobj
8 0 obj
<</Type/ExtGState/BM/Normal/CA 1>>
endobj
9 0 obj
<</Type/Font/Subtype/TrueType/Name/F2/BaseFont/BCDFEE+Calibri/Encoding/WinAnsiEncoding/FontDescriptor 10 0 R/FirstChar 32/LastChar 122/Widths 221 0 R>>
endobj
10 0 obj
<</Type/FontDescriptor/FontName/BCDFEE+Calibri/Flags 32/ItalicAngle 0/Ascent 750/Descent -250/CapHeight 750/AvgWidth 521/MaxWidth 1743/FontWeight 400/XHeight 250/StemV 52/FontBBox[ -503 -250 1240 750] /FontFile2 222 0 R>>
endobj
11 0 obj
<</Type/Page/Parent 2 0 R/Resources<</Font<</F2 9 0 R>>/ExtGState<</GS7 7 0 R/GS8 8 0 R>>/ProcSet[/PDF/Text/ImageB/ImageC/ImageI] >>/MediaBox[ 0 0 612 792] /Contents 12 0 R/Group<</Type/Group/S/Transparency/CS/DeviceRGB>>/Tabs/S/StructParents 1>>
endobj
12 0 obj
<</Filter/FlateDecode/Length 2405>>
stream
x��[�n�F}7��G����/AQ�M�4E��������P��Z�T��ҿ�̬(9�6ZD� �)�\��̙���lٷ�^�z��K.~)������w߱�=e���$<���,a)�f�d]}z��7�==������GɄ��fW���%L�,��,	�Rvu罸��Mk�z��߽8=ap-3vU���8��]�|z�V��|��)c������%���G$C#�%Wډ����X$Qk�YT-b��)�?׀a���0<c������\E���D���:��BD�r�ñ��,8�g���Vb�2*�@�����8,����5��ũ���[xCִ�N��L��������W{�6^��o��c�]�؄qnO�#8eW ��ޯZF����>���y�E�Ѵ��zv�����5�A����&]_�6Oٳj�����
��
5B��m��X.�{Ж�*������oB�x	�!2׏�PG��i�B��V�Tɐ@�Y4E�f5�A�uuߡL��b��U��Z!(�\�"賞L�E�;c�K��nc�v��"�B�@g)�顔�X6���G�ȳ�1��A���f�/9�3�2�D�Z/�5���KT�b:�'p`59�/-�K��q�g�lGUנe���b��` ��^w��%� ��oCn��[~��&�5S�+���4�Wı"�T�]��m}�⟠��C��[kJE�n��E(�"ZX�,� 
�ڣJe�k�)4�^CLb#����8�s�Hr�.8}D�aע3�Ng.Pt<���S '��e�38�$�&w��]pIv�@TD��&^���yD�"89
-AŇH.8+m�tBZA"㑇'�f�8@N2���T.Do�o@RB�k�	��� ���� ���)���*���d0���&�h��X�S��(��@'%f�������b��J
�n�\@�S$O������a.p=œ޾���~!g-B4N�����X+�V>�Uf���Prr���	����_�gl�w(kHuq3x����e"�,\?�Rp����pA"��h0���n�ȂW+|���n�,�|��_q�p|�~p~T�s�ȃ�㸽���9"� &�s*f�������W�SdX؍�C�*<w����ф2c����C9�m~ ��#�j:@�G�Tɍ�͵$ۺ�K�E��S��_�U�"_��r,"�F��LQ�%8Ӝ�(9�~[��𠪧��w7�<93�0�_
_�����j�E���>���;����:^�H�Up24�t����s�蘱&#vo�/yf�B��k���\���0�g�*#�����W�����|��u	Oh�j�ԴO#�٠�S^e���ėM��~\v�o�\�g�G	G��2��D��{@
�e&�*sA�7�_��1��߳��n�/�4nYV���	�nL�g�.蛡��`��5�!�o���N�I!g����1��F 7��F�X��R�$�8H���g%�$�Z7�)y�Ć<�|ݯ�D�=��i�}��vm;mzH�;���Њ�
���ң%��'�iJ��n�h%|��<9ұ��:7;�%���c�CM�W��τ6{r@���9BBG�z���3dTa�	ω�)�	�Gr��c��.H+����G��g;i�:h����`�N��+�R)���`�TMH.�!2����:������#`><��h'X�'�q�qAz�~ok�p��4�"Ƃ���ـj1N��%�C��}f.L��a�*\?�#�N�Ӊ9O��ඥB��Yp�ĉ�GX�D����0O�U0����ӈ�4�� ��4��{�.�a�Up�Ѕ��ap��E��p�N*+}��48Y�����d�-�Hծ��ƂUW�j_�%��$�t��`>���S��F���O���Z	QL�$��(
�z��1TP�E1ۮ,R5`6݄�66���>�=�v>X�F=�`{�.��*(�}mƚHg|��:ҙG�,�K��9DI����>na����Sb8?"�S����jUl�<^X�� ��[6�Xf�m0(��1�3�������z|:��Y���p�s���ٻ�"N�O�+t�a'+����͌�~����\ ��VN��V;+dU9��ܱ��A�H��|��v�x�	�EW�#`�n�z��<�cJE��\�nu�SZHX���]?��j�w��xj�Z��8D��5"Q.H{��f��<����v�s�|[7œ����sv5���&�n��û��b�$s	�#���g��:h��0�y@�(�-���]�i  �-;T@=��#�$;N`F)���,��`�0�H�D�}t�L�)l�v�9�m3uJS������bd�m�:�㾢��O�G�-?B_+�ڸ~�.5�	c�.
endstream
endobj
13 0 obj
<</Author(BiServ) /Creator(�� M i c r o s o f t �   W o r d   2 0 1 6) /CreationDate(D:20260107152052+01'00') /ModDate(D:20260107152052+01'00') /Producer(�� M i c r o s o f t �   W o r d   2 0 1 6) >>
endobj
22 0 obj
<</Type/ObjStm/N 204/First 1787/Filter/FlateDecode/Length 2768>>
stream
x��[M�7���q���7	�| �l�c`F�Xk2#cH���"K�h̒��sX����+V�{d���&3�M
�Vc]1.b��������⌫&�d�d��p�Č��$�����LN�%���.�Rq���&l�j2��r����ӱ�.x�ےa���	��hq�v�L& /�h��f�$�]��D�	�S'�]��荛���ф��c�"�t���pߣ.� {1c��EKA�����)j.�^^�=�r%��*�`�Võ	�g
��-�M8F�2B�)���G?p��\���[�#S��|^�=��gjO�A{��)��*:](��dA�&���P�B�[j��p)x��e��a����Gث��΀!�3x~�T(��RX�\�w�]�	A���`rDd'~�螈��R�Rd'4�9�
v
5G�eI���HX�9���`ѼZ0��28wlB*��Z��!�!�D7�I~��H�G�C� X�G��))R������"׎؛���7���ت���Z2���'dG����BbI5٥��7�ॅvrh����.�����)�ɹ�ȅ�}��gs%��L��E ʔIiء#��f�+�:�T�u(��fJ�dZ*�RI<���rNt3 ��\*�\H��U'���:�?6� (���:�R�uȪ6뉨E�!�ڬCY� �X9�X�L�L-� �T+��z��u1�([�R<9�Kn��Đ��Sfrc&��"����i삮@EJw!*���",�t^�B6
�cy+��X7��*�:i�S��Q��
���=�9���YBm��xa���4�a/G�#��(H6
������;H&hT'��D}���}�$귑2���(�<PZ�\hWI�]-�׮6ޓʞ�d�6u���ܸB6,٨��#�����8I�Fb��'i9�o}!_|�%)P_�)�
a`v"J�8�q�ō�oi4�6�42�_}�yI��d^mn67����?>�67��O����w�o�������l~zc�_���;���_�����/���g��������glF�1"�5�V���{����<�|X�>�l�V��+ۗ�����vH���N�&2z�l�7�o|߄���|��ӡT4 ��sw��(F��X4 C�\v ��+9�|�C�i �r��@gR�q���\5 C�^q u��@�m��X ��u'Ɂh���X�@ı�IQ���b��X�@ı��Q�����E�X ��g�X%�4��P��"N}vKNt��d�X0�`�B���,�:�S�8*����jR�@����Y��A�5y�~��yjY0㕞w"d�0�����E����	Ck �Ĺs���+�9�c�`�P�L\ę�̟H�P����5 d[��W��WD*��"� ,q�T�"��IC+ ��%�Ej�b�X�!�����IU|(���0C-k �b��@(��C!U#fw`<�k��*(�PD'�Ϧq�h�AX e��t'��*<��0��i���*՝_�P-jvƳ�a���~֜��������x�� ,�5U���+����s�Gd�]��V#�1@&d�m�s�{2�>Gt�iw5B\��V#�%�u�#�Tu<�x!�����.�@W.x�x�,HO!hO!��r(�(a�*a��C��O�VбB�����A5�A�A�A�AjAk
'(E!(E!(E!�[���<ty��<Ou\���ux�檐��^�i�hD}�;nAAAA��8\������8���	�S@xAqAqAqAqAq���YǑu̕.��7��$����#pR�x��������4�4�4�4�f��3KbFr��r��r��&fdbF�*31��j j ���<9ga�B�x�.(K!(Kei ei ei ei ei $�+ $�+ �k ֳ3�ggZ�δ��i=;�zv���L�ֳٙ3-�y��<Qe��2OT\<�����\���'��W*-�*ma��x\���*�qa�VƫO^?������i �) ��7��7��7Ģ7ҕ�P�\³��׾a�[��������cE� E_Y�����nR{<&� �c�
b� �XA�2V�
b� �XA*���T�����ߙ���bs�u���P߲.zi�}$��*�%�>4K�L����q�br���;�~z��ぱ�pX���d~��o.�E%�a�/�x�0/�奬���1�jB^��+�x�/��K������"s�y��%�����}��J��Bܩtu*ܜ
�çW��F���ߞ����u�OL?e��a�׏�ݫ��yu�����`���r��d�U�4i�S���b�����1����������ۿ^��_�onv��͏����cߧ6���������[�!��f�����������iG�9<������_��3��vG��q��������������ww��û''n��޲�vo��m�����}z�+w����G����@V��߾?<v��[+ɋO���'�}��4/���o����ο&[�i��w6���r�9���	���W͟/A?_�}ii��:_^u{�������<_�8\�w���|A����R�W=_��|-��e%��Р�^Ymp�f���,�`��2���ϵ���W�k_Jo����i���?C������_~�?���.
endstream
endobj
219 0 obj
[ 226 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 276 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 532 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 418 0 503 0 0 0 0 255 0 0 0 0 538 0 0 355 0 347] 
endobj
220 0 obj
<</Filter/FlateDecode/Length 21336/Length1 82488>>
stream
x��\�U���y߹߇� 3�3��w�	# �`
4-�,�nj�Y�e�-ݶ���)����ni�e��]�����=�}D˾�ow��������9����9�9g��B	!:��HSEYy��K_�j�Ҋ�)�^����P����iu�����|N]��Z7w�}�����#�oj9��Z�P�aB���]�y���}\v?!�%D~���-�|NM��݄X�jokn���.��T�^^;ԻL/B�҉틻�_������;Z�oܱ:���O[ܼ�3�.ã��孋ۺ�o�xӹ�&B�\zN�⶷�^� �0</�Ύ��#Y�a��ή��o�O/%d����w	��ݳO㮜�-����X9���3�R�l�w��*beӡ��p�I�0����{��jE������Y��H/ё4��]���7�s)�E��n"&2�M�lh2�?O∌pZ)ǋD<':D��=$�|hV�ڮ��Z	�Ǿ� ��s@,��#ְ����xo�s���H�ɺV[��^[���?Cf��]t�Sc˭?1��n��+'��׉�y&?t�-��獛?���g�'�H<?�/�`���Ԍ�����_ٯ�K�)o0�g�'����d_^%��zO�/}�������|�KR�=E
OΣ�^�A�/I��=���#�m/C���$$?G�[����[H~���K6��:��@���y�vB���$$�\D����g�L���sG�߇$$!	IHB���$$!	IHB�Kd���	}�IHB���$$!	IHB���$$!��zӯ݃��$$!	IHB���$$!	IHB���$$!	IHB���$$!	IHB���$$!	IHB���$$!	IHB�����{�������OR��qۈ���Db�;ܩI)$�d:i#�H�"�d7�\`.��������R�`��S���/����D
�TCc�#���d�'k�ޞ�5�øS����o�:�G$��`�����i.�߳8��B����\7ڑ�V�r����G5��oCt�p�������������Kw弹sΘ=���[_7s��iSk��TWy&WV�O*��.-�P\TX�?>/��LOKv�m	���N�V*�2�D,�9J�*l�MV���'r�<�t��5��y���gS�e|�&���Ēn(�ऒn,�-Iu�bR��f��Y}�m�:kFܯ+�5Z}��}�p/r	5$�㡆�"����M�
_��}M��^�R1�6�M��F�J�U/���O�K�p�%W�sD�f������V������F�F&	m�$�|R�-�B�gr��?mOߕ:2�)U�jkm>���7C�>���o�O��K���RV��!���l��T4V3s��'��l־/	t�6x�DKs�"��$�q�M�?rO�o�C_|<��n2������F?q�R}\��3��e9�#9�՛l�,TM��sۣ}���i�}��ߐo���-��m}��r�[}��]7���X+�3\P��	���aF��e��E�ʰ �,��*�j��I>����sU��~Y+��ʱ��-ی��$;�N�ո5��F�_�$�����u���dl�����`����}����F%�Η�<.^x�P�vR��l�R�����F-0X+�b++��KH���[�����K��ځo��aY<�:�c�o�G��.�}�}�1m��0�'|�)���Y�R�m�c:xB��`���x?9��������3������&�h��L�6��l�6�C��ll��B|k�l53f5�Β�R���)���7	�`e�q$�Bz��MzNʮɶ��l5u}�q[�Ab�7-qT5_���f%�n��f�Ug��k����w��:+��Y���>[]C�Q��̆���Qa���ԗ����S�o�kg���ںY;u�௭o�s���T�؟y;apV�Y��%�,�Z�		�P޸�MH��+B�e��&�Q�2��M7b��&B�[�1� E���a������\������^.��oꣶ��l%����|
[[�Oi+c�Rf/E��٥01h�5����L�b�8y֤u �o�?`l���v��<�~���Mf��ɾޖf��m`u����F��#B�*�Z�[��B6�R�(����ט�ڰ�Q��:��
!�ئ���j��e	�&�

�9��5��IxX#:I����� ���
���:�긖*�hi�%Q�hTaf6,ޮT+|r'4��^�d���.ml���5��l�O	=r�qe�x��X_�{t�}�53c�̴-���uZhI
�>������-�����`��*e#W��y{�@�n�y�c$=��661�q'Ll��w��7;5=Mv�U-���d������G	F��L4�`���z�An刈w�V�nЃ�">�G�O2��Ϸ$>
�;@���=`�%U�nL�ʉ-|1�狈�/ ��y�\`0h& �V�%�<{�bW~�A�l�|&�儻�`�(��D�I��(�N�2h���:Ѓ�GAe��h1�H��J[��Z�B+԰	��?�l��ǥ��ǥ�B|�8�y����G�!>Œ���h��1�#ć��#��8䏓���_���a�w����~���M�_o`��1��U�+��/!"^D���3�y�s�g��� ����	K���I��}�����!� �6A<��݈]��;����[~D�ߔ�!��Mـ? @܏،��o�܋��ݍ�q'����c��!6!6"nC܊�-6}�f�~�7�7 ��z�!6 �E\���q6��_��ч��+�A�F\��q	�b�1p��
q!b%���������"z݈��.�D'���8�q6�,�"�BD;�L�D�т��hF4!�!�"� �@�F�B4�c��#NCx��:�L��t�4�TD-b
�Q��Bx���
D9b�1�F�"Jň"D!��] �G�G�!r9�lD"�!���h'�\ht"�i�T�8D
"��p �~C a�؄N�
�h�",�8�aB��D4�BD�"�	�hC�:��A�*��@ȱMB�F	B�!x��"�È!������"�A|-<�~%��~�ƣ��#�@|�8���)bq�	�c�G�����G� C�G���!�����x�5	�?���M�_�Q�7�Q����!^Ŧ_A������D��x�3�{��Y��~�3X�il�O�?b�B<��{�U؇���^?���A<�x�0b7b�!lz'6=�M����#Dl�mE���Xb�������!��GºK��GN܍��Y��9p�?r���ș����n���&,��܆Enż�b�[0u3��	��p#��t��X�:�ĵإk���Xr=�*��:,y%�
D�?�p�?���q`�?b`�?�p�?b6�R̻K^�E.ro�VX>�x,都Z}t���,~�~P��?�> z?�f��@���nл@��������t�F��햛Ao�荠7�^z��kA��Z�nYz�:�+A'ʹ�c�4b��]�g���06��K�z6��K���9�ň�g!!�E~C!� ����C�"rو,����LD"�G�Z���CP�
�D(r�!��Y�%���OAA�~�1�GηA�}�/�o�����U�W@}t7�.Ї@o�P�t����W��lʟ��Y�X�8у��(C?LD����r$"ΰ��y�������;���y�}9Q�Q��=���������ELA� �Ub2�Q�(G$ ��V��0#L#"���aQ�[�C�߃~z�[�7�_�~�%�QпCT� ����A�z�=п���= ��ЧA��GЧ@�}t�^�����n�
z�>7�>^�� �Я��mG��nY�hC�"Z�͈&�<�\���وY�FD�t�i/��B8���4D*b"��HB8v�M"#D�!(���};0 :�!8�eЗ@����A�}�Yp�N��x��R�i��:-{z�m�����^�y�W��he�J^��8��o��\�Y�=�
�hE�
Nq�g�w��e^�2�:����9�s�����i��� �w�l�������z�*{{���" �#=T���=JMe��˻ts�Wԕ����tQ.��N�j���֮��JV:�+*�Rו����x:���;��:::Vul�x�C��c}��8w�\]y�g���Ŕ��D���yE�.n�P�7�г����gz�7��]�l��mn��8�{��M�y�9޹��x�p����<���l��Os�{���u�ޙ�gx�9�z����Y㝲��[��x�6{��=t���[��Y`!q���w$N�l2w��N�;�#f��t�ĭ2Rm�����.^b,1�c6�l�k�^���u�{�\�ޭ^��^D����v�v�v�������LЊ�h�ͣ��4�4�<M���jX�׹5��J�ڢvOv��b��T=MͯWS�ڙU�V'&U�������*�V9R*?S�[��r. ���VJ�/����Al��HK%�0e��J�&��5����l�l]�ױ�{�,�d��xg�n����~�M��E�����֭#������o�d.k����{�[��{ES�.�Y��;ui*\@�.Kw|�p�t������BX��=B��=�z�� �R��Rs�"�j��*�ɿC�����B`"�Y�t�Dd�����ys�?��F���1p|��l&���c�i�"�;U�&ry��G>&_��ཕ�Hj�)��?�8Q�//&j~�!�c����|˃f�e�"�qK ,0x�mx����%�	uu�3`=BǸR��4���5�Ho�2���t�.�C����
r>YI.$��%d5YC֒�����
r%YG�"����r-�@�#דȍ�7�&r3��x+��l��m�u���rn'w�{���ߓ;ȝ�nr����O� 6�`��l"��]`e��m|�H?�d��#���l';�;!���n�0y�"��`c����K�u/�G� O���ɟ`f<C���Y��/�yb��Rϓ?�`�$/���+�5�y��M�!�Yw���B�ס̛�R�B������ ��rX�/B�B��;���/)G�#�cѻA��MBY�Xt�����,Bw�����O�b�7��(��ߏ{��`t�߻���9��S�H�v������=>��q��_㝿�������g�{�{�{��!(ü��8ѷ���}V����ay�C�#X��?"�	�`���`� ��|F��G�簞����W`9�ZO�|_ߐo�1���dhLj褜!21��(O����
*�b*�5MF�TAUTM5T��I9���rT?�',a4�F�zi��4�a�4�8j��4aL^�h�rl4�ڃyQB͘Ѻ(aS6�f�epM�N��L�Cs�xZ �tHgA��2���d>9����#`U������>I6�	��>���N��~��� R�P7�$�K�w��	��œ�E��if�(Q����+�B.�S ^ʿ+6O���Ԓ��~7Q�[aY/��l+/��K�$G��"����qj��Ԗ+�����*�^�Փҡ��|.�
\�����uCO�\�32�>^/h���J%[���Mr�egg�p�9[��l9y�K��8����p,M�7���W%r���e�i��`	��xK�ڞm�����c�"��ˤIye6��g�I&sR�h6�k�}!�|w�����܇%����JN,�ݚ��i�P�֪��!�$��5�q�桛b���`�5�Y[�!�;�u�c�%�b�
;!{�JuF���R8��c��m��*�nv�ļ1*e�.�N��8�Mg�d����ΠcW5^��L�Ē<���$�$�P���YYY��up0K��c}�Wv�>;#���?�!���� �mTó�$jӏsX��8ͦ4v)Y�4g�3L*n�rQ�%#!!����)�\`7+���w�eXU4ZDԖ�|{�1)F���)$����R��X�S�L߽7j�(;Ok+��O�&j5P���.DA�CL$�\�q�O���6=1s���Do�Vj�;|��*��l��1��ܑ3T��cSa��2߂c�����z�.6�m'�'>+N$�q23��"���{�V�e%9��T��4�Y׽�>mx0��6���Ro���l�=K��[FG~��%5��[5��a�r�*a�f߬�'��"�K&��I�.�E�"Q4w��L�	��-p4l�+�4��L�g�K�{zpΠp��j��Ȅ�Ƽh��`��+Ǳn/�rs�gvn�ë=����N���oR�ej�*�pfAI�Ą䪶����$�T!��H�0����k��Y��UUC�)3��V���YN�uI]R�9F�¢��Q!�'È�$=J¹��:˭"rM3��V� ���IJK���E��4>�1�hn��g\����oť���«\U=�U���鬳�j\���_\���u$�/z����YC�i���_�'|:�$�L�M�V�[í�D;@5�u�pHb�OkխI�~	�	���؁��K�>��{'86>�������̅C���r�p+�e�"Z!��E"�F6��^&q�� �<�a2&���k���v�o���C�4�,��w�6���=@;��Y?��5��ddqVa}0IY*�ԛ�;�*���J�<�`5�$D*Tl�f�UtZ����$J�Za5؝�r�R��d�s���r�.�7���{���ĳ--2=)z�kt��.EzzB���n=I�mM�R�fG��]�.n'��W�0X��

��ZWPtkpI�}�G����paI���U3���~Q�_jM7i��W8�:.���ؒ�vZT���V[R�HJ�(��
>����Z�L%��n��OI�%$��
�ڴi��>]&*&�$����n��q�=DAbh�_� ���`N��c69a�y�D�M�{撋�X]Q�`�Z��ƒ��)J�ƒ֪�3�&.~���N)���.z��ڒK��<�wv��yTx/��?���]�c�������~����:B��D�X�U,V�#[U��l6�.�?��E�xq�#���q���%w.]3���6����<%��ݓ4�y�3|\̢����p�y��e?2֙�2gڢ��OՊ���:KI��@��a/+�I�}�2u���',�"=��S�~�J�
��Z[��#�� ��un^<>o�����hፔ��CT=�������9V_�1�]�����R߶��06wjN�8{�Ϋ�?�w�{Nv��p�B̋:�{����U��}ؑ���ɛ59W��K������=cʰEa�ao�F�#�K?p�n�Ҋtt�Vc�BOu�:�"#;�ѩ$,,Mz]@m�r$e����=_-�9�J.��O�~�h�&�)��p������|<�2�,��~�7��G�n����tbp#Ld���=D=$3�ǭT���4a�Lc�-q�ka��J=�
[N�A6����u���!<�HƼ;��	n[�v�x^,�.�>�y�Ƴ�OZ~����I�Qr1��;r<Y��c�k�sj�j9,w�X[���s��ֽzoo�&:.Jm�)t�L7^�9��nqX�q=%~Y��\H.�F�-��pgl󌟦��n�[�=!{|-�p��݊eS��y��x��y�rkWm6,ϖ��	�ESz�j�U
�Di�`l�����a��F8�鞄�s��DؒFV��H��"j��#{<L,��{|����"Opp�>Ɛ�~���s>��*��{�E��0�D!)�VgAܔs<	��b�o	��m�I��D�����2�3O���ظ]V�K��LL���.�5��Ӧ*����%s��r�42є��ר��i��]���ENzEZTTR�-�$Qk`q��Ď�S�؈^���|	[]j��ŋ�>�l�r��`�~>��܊��JeA�Q�7r�7@�����ab�@j�[S+�<��APص`iς���_��ؓw�dl��4�p��)����)q��eōg,Xט�=��y5+��q���cy-y��S#�R�sb3��	J�B$Rh�-�3���ڲ�՞	E��J�D�S�{2g���/���&�Of^��m�_�]$��赭���i�o�Rs`����i�i�1m���:Ƞ��D�qS���D�&�OĉD&8d���2��P�u�Q���4���ȣU�V�ߺM�w?�༹ptLe��9K��I�;���o��^�����_b�?�+�<!JR~{J�лƢ9�Z�2�r8Ppp�+��]�l��s�]ԹqA�Q~���ɮ�s�̙�n����DY���h��x�C+�=zYeYϦ��E�%N�s.����I<�$�2���عG��*�ж�����oM�TE��[���ظK_�gg�E���ƭ?]���g���p������u�U�T��*� )S�Ė�XG�Jeb�Ѭ
��/.���^ܘ�T���=J!����`R��*hƔ���)E��
�\�?	���Ƶ�����CGa�ft���~�7}��.����H$�����:����#��z�y/���ǄX�\[m�~l4�K�)%���C �f����?ub�8��;�/�-��̪+ͯ�3Fe֗���ҏ�v��.�p�ܮ��TO�pࢲ��Δi���)S;`g�0p��c�&�?S;�\�[Eb�
�¥�ռ��I�S+h�[�N�vh#�U��b���<���,F��o����ڌ9��lo�O�$�.x{������q�&����M�X����|�:��C�k��
�L�O,N:��.�A���udMthy�\��c7sW��I!�ǾC�W�[:��Y�:}d5Og��cV���c�d���-��A����ڗ�ǥj'I�m��Ý���~�*e��5�T;�Y�3/R�3�റ�x�^*QJ�+�\�0�a��I��;�S�#�Ű#<܎�T�c��X&z���9~�DsP��v��R��M�ErS��T�D��SԠIe�������k� �����`Vց,W)l��\�c�9�Y�1?��ǟx�����?��Lns�7�#��Ec\ �]���=FW��F)�ۛ^<I�w��*��^2�⣴jͩ���ȏy���{�����\��+{�?��g��n�"����x��.��L��nGX�'-�^i7��N�	?ݡ����#o܂+��9ˋe	�M��9)|\�=J)�������������]辿�[���6]�i)�(i���4	I�aE(���#���QDY������ �(�(��#��s�{IӲ3��������{߹�~�rϽ/�E�D$���r��'�y$7kP���/t�#U-�q�O�w� ��@OA�򪪻"���C8�9O�P������AY���P!S�WFzyG4��	/�OO�(�sm�ݴ���H�Lzg����Q������¿�9e��,}=�/~3<;"$!P*�ɍ�|���I��)t����:92��C�Zq!�=�cₓ�C�s�B���,�����ߢ�� 7�����|qd �wRo�����&>IM/��}-�=8}#<{?�zj�����3gaHH��������H�\,	��.J�Z�Te=zZ!��������^�S�ñB�q{|yIsUrB�fp@�AI�pN����̄�D�q���/'�NJn)	P\���n� ԟ}�8�΍4���(�����	�꼀���+�>^�a��P�B�2�ȑ)�#���5yQ��3�?!���F'q�E!�+��vf%&dd&�s�`��n�x<j7�K���V�}�$h����|��F���9�5�խ1��{�+[*�IC�����et^>��"�Z�Pf)-��Q$��ˢ�A�C�����:��9@~�R���Q��'�,X�7~z��_���0�_�t���0�ǐ��]�G~��K�B��[.��ǆ���K�S�(��بAa�B.�{#8>�<Ѡ��=B)��P*��y�+�yB� ��b����[�UD:��JDG�#�^P�#��낤�|��2�;��
<�����.E"��g�-�N�Z�1o��Qq>SFz�=<F��cC�b��=�i���󅰐�¢�b!_����nJ�<��Ó#������A�{��FH$"v��E�qyUʏ)������q��}��;qxF�9)	J�@���Ed%$dF�������J.�r�#���-w��W.�}�T&�FyzF�&&������x��)�	c��5ۚW�^I��@ 4��sЉ�{ ��%�TdR�8X����&��g��eD��q��2�^,GG���@��x\ˌM�<<��ظL��	Ⱥz&wr_�'А-��Ύ���2�g	1�؈cp�p~s��H;=�s�#e2��c`�럔�����<$��+f������cpRR��C�j��8�[Q��)�����+�*�(KG����=��8� r�����C�}�f,DAQ�I�Q��'"Hԙ��}ıs�o8vӞ��}~~�QOL�M�UB@��T"�A��8���0����ɑ��Fc�1��chG�Ů�SSt1:QI���Y�+��3}3�v]Yaffa���a���:��R�2j�̢��SM٦��w��=H]�_�2\0\���P��4�];\�^{�if�0��.*�H=�z�; N:�ǝc�#шA����訬̌�x�Ӈ�`?ׅ�?^��o���>��I/FoW2�2�bד���ii5z��:8s���7љ��1dZffy]왌ޯ �ň�.�7Z=fd�����Z��^x#���f]/�)���P�P��oа�2�L%0��D�(/��#u��l�����u"�9REP��H�.���E~��?R�ɕ������Õ���#22Fd@�p�����8��eys��&.��Ͷ��.O.xQ1�Yq{���I��ⲳc�������ψ�Bb��	Q����ޞ����<=9����Q�R���5�1(:@�V)k��(��!�E~Jȉ@��H	!���&|��NN!A�o������?�j���.�)iL[EV������9I�#�)}�iy��F4�&���vFDx��5����ş�Dw�;�9E�4�K�� ��:��Y�Yt�.J�����"5wD���S�BX���'n�Mh]?����+�t�F�K�4Z՟�a K_�7�h�hŝ�Xv[Zxk�P��w���H���� �]NZ���|������G���G���nr��m��o�"L���&7��Mnr�?���5�Mnr����&7��Mnr����&7��Mnr����&7��Mnr����&7��M�%T�&7��K���R8Q���x�.�{?�B<��N�<�P�6�<����|�?cy𿱼�h�{���H�?��b�.ay	��9������2"I$cy��@����h�a�_�)���$!(dy�\��\" p1��Y�*��������B"/pˋ?��^�=,/!��sI�� ��~A�Y^.�U�����a�'p��sY��3�3~fx������?3<�g�g�������3�3~fx����������g��<A�M����BKX	3a��z�}�Y	~�@�8��+���"���@4�5n��S�-�I9Q\��V��mz�QC�c�"�@s;�m�3�k�H(�1�L;�u�A91�Dpq�V���k@�d)�W� Zb+;Z�Ћ�6>�Ӟ�7`���S��@�����kԫ�^�o#���ZJ�Y�����n+���f��a�Q�߈�ʉR���c��Lدyx�K�&�yY��)�C���6S`qD��t�(0�^(���%��i�B���bcm �H�䐮vh�g�q��}u�1&+��� ����vl3�	[��HMx�S)�J=��|l��a�z6l��
hհ��"fa��4�#���Ei��&<+�ӆ=Շ �h��0k��[�gʄF6s�&����v�2�X;��3Gk���K�!v�y��c��m%^��ь�ښ��v�fv���ۑ}&6���L\�89�ǱF�kqZ�`l`elК�j��L�Z�Q��A+���]�ʣ$<���_y�
5�;��4C[GԲY���lАU��|�S���o�8t8;�iθ���kg���4�f&L ����?S�%�*���
�-��W^"{�"�qV�12;�aC�T �-�tC�(ٜK��P�"�v�� v����N#ƀ�c�L�ct�,Gm8�-�v��q(��L�iǞf<cwF�!�Z������>@r6+\k�����F��mk�:��Uƀ-d��a�(��������z��;��N��>��;�>�y�yZ�T�V�'-^O7�Y+k��4#^S�ʿ��h��$�|b���vÿ�[������g�q���΁��q�� ����9A8j��y���؄�斖2���UL=0��Uߌ�S�txo3���у$����:G�*nb#ӧݱB.'�F\���QU��z�gmp�:^��
�u���5��\		���V|�0�裨j�y�$�RY��������}'�ew��݀
��̡�
sf�T�c�����bdw�������[�r(rUΕcs9�0�f�@���Tlw����>�ssVj`���c&�,�9������l�#S4D�.?���	�pzH�mG~3��^ǮU-{�6a��{���m87Y���-����y�v���t.w����}w:�W7ŀ������F|�``�W��o���D�*��3s��.b��dF�o�.;,��cѳ;U�3�����a*q^%F'Ǻ�Kw�U����u���}�h�~l�7�����'��~Gs��e*Hh]��m�1S�u�ǎ7�_gNc-��٩ۄ��.�z���'nVS����Z�Ī����{���:���,5a��*��n��� ��VB���J�Z�`�T�R裠���J-�
��z�A����#5�C% 7�q�5�W@{�qE�ۨu�W�.4VE��s�@[5�Tc���[�*V�(����F|1���|0���(e�Di�SN��*�3:��CK�Kث����C���E��p�,b��c!�Hg *�-�;>�@�ϟ�mf�V`��:c�
#@3+Y[9�Z�
��W�gU>�A	F�����H1\��;D%�,ĖVc�X�!k�p��*&R��U�B�����;5~g��]����8|�O��/�}/����-&�U�c��*�X��g�3Q������)��ˠwd'3G�f>[W,���n�F-��c�H����|����9�4��|�J��r�r��j����T��j1[5v�٤��FJmhh��(�ަ���uJy��Ϊo�*-zSM�EO�i���v�hn0h)���nE#(��Π��G��Rk��F�DcҚ�Ӡw���D�4�lh��F��2��7[�Q�:�A�1R� c�I)��٪�Sn�ƪ��M:���7����̠՛l�<ʦ�S��:�N��QF����mZ�����s��v��hSh��:�͡��̠�јl��j���5Mc;�j�7R��:�QOY�0��� �@Ԯo��&8�j�[mJ��N��5�f��FY�`��shm
�֤�j5�ѐ�f��`���&�$mz;V`�,V3D��F���j�R�&�Fk�&ʎ|�`�h����T��+f&����0�0M��X3�mT���Ni�!�n�>8٪[��^�D5[�4��zl� n7�A-�$hb�Bɣm�X�ުt&�ǜ�(�QW�A��V�g��)�����V�Nߤ�NC��:���nA�Z3��d�۔e���-"I[�f{��n�IMՙ�6e�c����-����؞���\C� il�jl�f8��&�5[,F$���&���k�T3��%,�F��Bx�z�3�,��LP-V\Ղ�>5J���`����vl�#%�]�;f���G3(n�rA׬�+PJ��X� b��h�6� k�I&�����ْ`Hd���8h�Zf%A�C�mv�A�$�c��]y�	��*'V�zt�V�Ѭ�����qd��CL���@�Gf"�F���ߣP� q^+��:��(y@�7�� ��VPu`5�����6�&e�a����4J��!�RA���$BxqZ�u��ܼެ��`%ʐ�{��S�`r�'#7������_��˫Pplx!���=�����T�
Z"��f�c�D�S�:(x&�.֎<�s+ ��f�4(?`�A�2�5LM5�3	Hc?k�j�Z����pEd�pS9\kQ�K�)�tC����Sfn����V0^D�B��z����4�A�F�`Au]3Z�6��f	X�
����L�-���*��aJfѰ�� Z�M��-�f�	����(�2U��;�/�!�u���0)e�E���v�d��n`�1�)�%[#����V���P+��f�d2@�������[����,���VQ��T�����PUH��WC;^A�+�)�[C��:��fUYD�WL��*�(TP��UjUu5U��J˫�JU�WZQP6������**ao/��Jk*)4!��TU�����%��UZVZ3AA��T �E�4���Wה�-�WSUc�U��*���V�V�aU�����
�T�Р�K����T�c��+����.-.��J*�
U�9J��G����������rU�_�_�£*A����ƕ�p̗�ԔVV 3
*+j��T�����q��*��.�F)RW�z�NQ����
����A�ժ>,���2�U��
+��G�G��oݏ��G��~<��� =�#�#�#�#��������c�w܏
܏
܏
����d�� z����^�7�	2>K�o���U�]*�� CZ�T^.��;�T���c`w$���K�T���?v��>> ������
�}�GzQd0�B�CH�"�#ƒ��)�
bw4��G̅я���z����<�SzjA��AO;�y F���X�_��' �Ă�4�3�����A�T��z悞'a�*��0@�i=A�'�d��B�Sz�@�	�� =��e0�Y���_g���ГzrAO)�=��z怞'@�Z�H�诇;�EO�Q������L=�3�,==�`�.�>��G$&D�����2�Y�g�$�"��S�N]�����L�����Sm>!XN]��n�r{��)S�)̫��/��Kxg��n!�WțrI�")��^f�.p�r������%�"���Hx��ѣW���P&�u���!�����q.��������G��SX`b)f�9��Xd|B, ��RR,?���}�'@���$�b�	��P`9�!�D@JDtG;�R(׺��ɹ��ׇ:�"�B)d!v�av�xK�J8����D)�B�x����%2R�q�r^mFt�>N�$�񵞷�z��U؆@_m�
I�X �|��As�^���l�PH
�X��r��* �l[��CJXoV��J���l����m�qv[vl��ebL}p�q�]��ݽ�Z�LH�� b��!L=�o�tx�z�<�&h���Y�uZ�'E ��N	��8Pl�#t����-øe���l����C/=e<eD�;���}�}2���I��ܷ� �Hn�9`�u��E�\W������w��<��K��<�������{�ze|W� �)�3����X���-E�t �9y�������r���R�����M,��1|-��:�om2)��v�QA����ޭz���U����5i���8�'�]_R�R�3�I�8i~��+rR����]�8$�&��~���'h�@�, ydg��uU�ch�KO��Y��PL���o�w��>q8":�EϷ�g��/�MzVsjމ�'���4vWWg�X����������O�ȁC7|Ƚ��Nx-w�%������	|8c��|ho��H�il�S��lJ�=P��G����&]Z8�z$>~7�5��H:]���]�14�S��&UU�O��Ӳ��tNZNVnf�Dh�4��[�drZ��K}x�U�x:�i��
�h��ZE��+����R2rr�SF�E9i�t4cQ�M-�fӝd���I>��$=	�p:��r�[�V����ky�߈�m�����'�o�_�7g����e�=�O�Mۯj��g��+[�c�$���.�<o��	���z�����w�ut����Gi}-�xYx���<���WiI��?|x&�����>������X��&��]3�?�yi�K�%���	CM}:d��S�6Z�ް���!/�qx��5���$�{$b��I1&����8�sn|�1E����F�|�n���wO�'��4fFm�䯿�9����Q/�y�<hwFWg�I:[>·CEv\z%����ޟ�͹��}.�����<§���a<���o̘w�x���.�2,�a�´�N�CaѼ@��ot�Տ�E��#�h�ck��}Y[=�$�+��K���T��g�Z�q�/"X�Po*�Hߖ�#�""d�D��,L>_H��2z4]�hӜ�C�	Z[[o6��z�v����h�C%W4`ArQ�DkW+�Ƭ~[�3n�u����N-��~�ٲWR�7~�0��値_����m{k��M�Ox>P�w�kSt`[]^�`������y�􎦏�G��Fl:P���j��US>�nz����%3gf��!xS��wĨz�>&��۪�N�@4�^.��(�Ƕx��5��-�u�J�p��[pׇ�)Ou��[y�Z���z՞�����w]�ǹO~��1{Ib�s�Ѽ�.��~�Ө��!
zU�������vR��ם{�Y9���ʖ`��_�T���Mw
H(cߺ����.�:cvշ����w�����?�X$�q̢�p���SՆ�@�~�+W�:7--��d�Y_���)����[\������;b�	]1���Zܔk���e���m_{��C2�᏷�����Nrی#������;�������Iz�L�jv >𫄈_y������{�Y��Zj�y7��t�����ˎ��}�����ڵ��h�}�����y�Nܵ�ħ�w����l���=�El�[�Ɓ�[�t���j������'��8}ڑ�E-��^cJ���8TR�V��������z��~=��3�����{��0�����>Od,�,I��f���׫�1%N�})�4��]}��9��,�HSnbQ�q��e"ҹR�.���ɺ�ǧ�������v��}��2Z�.{�=[L��4�t:j�}��3h:-=Y�Kg�e�5)���2S2�3rSr3��St�Yi������zm�Xb�}U���o99Qۚ6n�<u�x�
e��p�t�<�,�F�{zK�sR�\\5.%p,�����8��m���2n�{y8G�_��NI�#>�fա��5c�>����c{>����������?r�k�'=u�wnB7_�svE����_�d�w���ۇE��7m��#1q��G�O��"��~~����œ~M�|hգ�s�U��u��ةN��.o�:�h�s�:z�>l�pe�8n�^Ӝ���^ٚZU���E�´�m�/OΈ�LZ�Z�>g����J[��l�:��+�ߘ��&��dóN[�`�q��{TG�*fo�	.~dٺ�nS�[W�#}O=/���;������0gu��MTϼz��X�-��w�����^����ؘ��m%�������#�>�]p��U�16�=pVE�yQd���_��+��V;���ѯ�>ҫ<��g���v|ˮi��1>`�ۅu�:|r�5��M�E_u�ٲq�ڝ�_R���Gם��tm��4���u9�)U#�>V�%}����;����g��?�船��n������n�8�t÷KZ�����u�-G�r���w�����?͚JV�2۶��IQ#��<���Kק~�а�߽�Y�x���e-��/�?����y���K�9ǹk`�&p��$��L\�Ca���T"~"n��?)td�?�1-���)v&+�a2S7c���l��	�k�7h5v=��lo4[�vT��:��HK�ʠCqOO��5�sg�V�W�6n9�I�IӔA�������DWm|�t`E��_����v���N�A�S~��CF=�i�d:�cb�7�@�yŃ���G2bX��/��k��0�������FW~����w�~��ͣxk~��dÇ	�Uo���W	E���W�U��qL}�1�������yr��o"�μz��g���&�+��V������7,=��`��5��]�]�+�\5���m=䊰*�<.�~�g�E���Ԭz)�-?����g��<�Z��&�r���/��D�U��;ߛ��Q�_ ���=��Os�å���t��w�'��7����=��D=={S�g?F�~x��ǋ�SF��/�*��Z���&�{v��Y͟���^��W��Z���6���ROW1�B)�PWAW��w~.v^F�ًJ9�j\6���.t�r��31����z��a��҅�&s�O����O�iSNnQڧOj�������>�C���5���v����|����1�q�^�"��0r����~z�݋y�_������/.W���|�s������_/�I�:����I1Q�?~�v�m�R~E��ew`��G�I�O�X=��)�x\��<��CԈ/���Mݒ6,�*=t�2�w���̛�#�?��]�C��J�{���O:������?Їw��'O"$�'>�]������oMI=����G��~�Ҳ�����k�o�3�/�y:1S�\������҃�]��~�����}��{֎�ӣŵH��M�XT�{�����V���9�?���Q��>�LT��&�뗒���O��*�K*��g��K�}�|��!�=����Z"�x�so|ͫ[�[��E�i��so���� ����Ɨ{Ό9�(���=+���Kyi£;�E~�m�a�+m5���U/.޼�텭]K��?z�����"SפE�ot]�{8��w�o�����Ro^ ����צ뗾����q`��S�!�O�#��ʱ����Y{��Π;�u����x+������R��i�Y��w� ���`��M��3�F6n�Ѩ��c��ܸwp���������V�U$ ���Fު&_�]��E(�w���~�j������<rwͳ�	���`qh&ۆ�WE�.w�V���MIP�Y?�s�ˌ�K�go��9���J�uU��O�<� ��2��Q�������7�l��qD��tu��ӹ��b�}q���"eM^�iŲ����&�x|���jL�RO�����b���c�(y�0�EUE���{��x��yb���M�m�7�6�ľ��o���P?��k�u�G���3����v���,�.�m���6Q�T��e^J}�9�k%�[N�����=�Å��=S��P,Q����vF]�Bu����������(/_��&Q>롆����G����킎l�Wa�p�*Z����X�@���?�Y�������WB��[.���Gb�K�듃���=W���m����d�o7����4X����������ݐ��������z?��\.��lymzó����M�-�����/����6��F�N�������.�G8}�^Y�_2�{ޏ
��؄�����[nm��7��˴{��̸��ZG��|�;_b���'�~�$\��C0xA�3�#j��Q)#�x�t��'8�a�{�j�qËʝ&Q��4���w�w�'I�>�|̵��
������8�j.� ����s"���c~�A�|��X�4N1h�$=f��f{�uL�bƄ�Y��6@�e�&U&�e��8�`20�3R�e�aHeH�����5�򊡫�R�k��d�u��?�-�� �RJ��t����&O��4��R%τ���z:v?]�m�����)���+μ��_�t���Ԗ	��n�7x&�\���l��ta����v�z����J/��U�|�壗)']l+��?�.�P������֡.��KV���~��+Co�-{���dy�̼�Ӟ49���M���{M�穮{�^�텻����Ԙ>×ϖ�G�5��F�>�==o��%�1�C�֮{���mю@��Bu���_��ӱRȜ�)�3#/�����l��4��}Ӹl�����^&_��uy�S��Ňc����&�Mo���Obg�?<�t��w�Ɏ����۱��]d�X*/�/1q�;ǤY��w<Χ��^������L��pm�����ӗrz{�l����yt�����r��.-Z4��J��T�տݕ����?{���G�K+�޼2�Y)����f��g���~���*�z���,>}���&O��87��C���
A#Ū��\��8�$����a~��N�.��j���[9����ܬ�A�¼Ug�X64��abd4h�:���@��Ȃ�#����9�y�g^��@���eE�Y�Eی3i�3�]W��n�m���a�$-<�a!�4�.Q�<9h�Z�
Μ�-��V7�412�-�8����r����I�k�
��;�[���%k�?7���f����kOq��(�뛲�ΎX�ՋݏZ�.�����o���*�P;��++َO�N��V�PX�bbȼR)|G�ѭ���^G߽���;d��r㝗�Nn��O��>�;��|�^�����O��l|�K+�M��Z}�E�krH���@��a2�oL�������,��Ud_�x��FM���ZͿN��X�f�}��˯�
=��?e]��3\��/o�֔~2����+3�.lb� 6OTq�f��$
';�c�iCJ���I�1c��.�j�863452�(�i�P�7�w��Z�[��u�.w,XѺL��"z)�ئ�Mf�[Q~)��A����jw�Yqb��cn����U�F+�/]��l�|��]�o�)ţ���&:�<��l09�������[u�����Qg��Oe�]�MKNn���h��}C�0K��%��n0rx��W������L'/K��Y���k�8=�С��̭��d��=Bs���BKO{d��������ً޳�\8=7�N�n�����2�E�o��N���]x��ƫ+����K�X����Vc���ُ5fy�jm�ͫ{c�տ��{�� m� 
endstream
endobj
221 0 obj
[ 226 0 0 0 0 0 0 0 303 303 0 0 250 306 252 386 0 507 507 507 507 0 0 0 0 0 268 0 0 0 0 463 0 579 0 533 615 488 459 631 623 252 0 0 420 855 646 662 517 0 543 459 487 642 567 890 519 487 0 0 0 0 0 0 0 479 525 423 525 498 305 471 525 230 239 455 230 799 525 527 525 525 349 391 335 525 452 715 433 453 395] 
endobj
222 0 obj
<</Filter/FlateDecode/Length 54751/Length1 144100>>
stream
x��}\T���;���R�*��.����]4FV�"���Y��K0V�XI��Ĕ��M�&YV��j�{o7���DS�MrsM���� ����~���/<�y杙��̙�3k � ".&�*�/,���j7��6����O+xm����O^�ж	�s����}DbjU�̯^x釮uDg\Nd�R�l�s��w�jB�������PJ�p/�5{v�Y�-ފ����M���s�kw��"o�8������Hw�3銩���
�/��nmXPS�Z�U=H\܀�S�W�X�ך9�sP�9�ni���lYFZ�V��;�z~ݍ��I��=D��,\�di��6�?�����u�f�w%Z���}Mr,B�R�u�#~�����׫_��v��	��?��ׂ{RiĆz!t�Ğ�-��߿%l���u�*=�^t3�h�i��H;�Ր����%d&���@��Ƭ�B4��m�4ͤk�Ϩo�n��hl�d���D����7j�N�2O�i��=�xSԡֈ��o&�f*��c�����i�����3��j���G���P}�tr����놼���:v��4��W�aJ?��=b���l�}�=��_3��v�S��gQ?��v����}���Lt��<�?f^�u��M���ێ�t��j8*ފC���ߎ��������r��c�	�}/=v��n�?��+ӟ�8�V���1��u*(�{n��N�~(-d$=����=���s����4�d��ѾAt�>�*����*C> �l�a������=�E�r-eXޤS�u=�2N�~Ȳ�+����!a�G����y�}�|�=(C�C���uD_�k�o���e��n�I|����L��c���k:�喝����| �����q�4*;V���{)�_P���p�1�2�8J-��~���e����S��@�涣����z�7Q�Q��Tq�X�V*�>�m��c�6-���U�K�+5�����A�A̠����@�Qu�O�~�/>%����'��-���Rm9����}�o5�k/�ޭZЂ46�:�������VE�-����X�wzP3�U���л��>"�Q�[�wp�q���Xy��M�+OT��:�.�w���L{�\�^���<G�ە�3��b`6�<n���U?���K�B�J��+�s�f��?���8���;^9�3�>*��Q��'>���
��_����k�h�VB}���:'QNkm/=ѽ�������ؿ�o�2�G��=�*�R�H���.���J�;袎�H��#��f#Uj�p�v��5Q�v:��x�O)�TD��J�.8��N���-hAZЂ��-h������L}�4�	>ge����ϛ�g���L���e?���-hAZЂ��-hAZЂv��q�=hAZЂ��-hAZЂ��-hA��L[HC� 8����ߺG=� &���k����hOЂ��-hAZЂ��-hAZЂ��-hAZЂ��-hD���-Z�~g�H�$%A
J�N&q��&3�@Y)�zR��G���&R��-tm�]��64�wj�����SG��;Ü6g�s�s��<�E/�bj7�R�8�����8tM�j#��#N�ԁ���3�#����͈C�#�D� �zT��;�5ړz�>���z㡯}Y�����O7}����ɿh�9K��C�&����=�-�R9z�X�*ݣ/ֽz�R�2������ETJ�S%�@�9�u΢�B��&�E7�CL�b��+��(��5�|q��P\"�;�n�xJ<-^0�&��Xd��b���"~2Z�ӑi-�7�4�m�F:M���:�U�Hߧ��ש��jɿ�FG�]ڡ�ӑ#pD3���8A�~o�;�ԃY>͓*���7�Ǻ$w��K�,^�p���Θ7w�����Y3gL�6����)�<�l���N+[2ftqQaA�(w��SG�2|X��!�s����#3��+ݑc��F��YBC�&]Ի�U\��eV�L��1c�ȴ���N�*�������UF1��%�(YDI7�tw�6�ѧ������X�r���2/��BW�ӷ���m�4V$��P�Y�4���U�"_�9�EU���^�*��ӛZ�# #�|=\[E���Z���Y��>=����7��[ThOK�0|T`���B�Xι��t�������l4�*;��U[=��ӫQ�Y/jn�����t�z��,	]���v��]V:���gΰ���?�ڷ�pOu��a����]�&�+MhZ����ɶ\��YH��ʼ�v�,���9�>�J��V9	�Ӥr:�W���*�
|/���k�����o|g��N��Y5�f���fWa!�[���.�pW�Z��/嫫Љ�rʼ��B_�+����`�d�Q%P�_࣪�@-_NQ�l������(c�ʼ�h`�ǭ���m�QU�v��P2�����>G����鵧���
���B>%����c�.͸�Q};��*,{�aqz5�^!��b\\�#�a��2���pz��T1�%PB��� �g��Y��Z0ƞV���M��d��Y:Ų���&��q�ƥe�z:��
;5��@ю�NM�E�ƨa��s���3�r���pɧ����D��U�pa�'ze��XϷt�����k<��,)?,�����Q�UB+�,ζ��j�G��#�KT�K�������9����*|�+\�Yٮ4��>�[-�V^U��Z���U\�������iVs��ݼ��j�p��fWIm�k�w��h�$��Jy�X*����Q~�Kl*ku�M�+��lD�M�^�&����������r�`x5�N�pʄ�4		�Q޾�M�d����id�,�'��Mc��o�i�ȍ�]M��sܪ�	>���t�@irl2���L�V��7�-�0w�f�0������-RX��1'�6����2"M
�lBI�k���X�@�w�s��J�HB|���0��`�}R䬕�ouŜ�
�{P"�*��O�F�Os�D�C"}ᮺ|_�+_��?��!���/��t��\؈�b�d��t����^�M{Ѿ�"kiP���e��f��r�%���k���� �W��(����TQ���a�(Qlԑ��j0ת]��[GS��"[��;��X�6�q��drLs��QNEs�k���`��gl����d/{�H�f<H��hy�Y5UN�#����engO�|Sf��p{ �d��k�/�/�[ꈾr�1g�VTp���@���@�2;e�FY%�-�ވ�ʢ��0em4ɵ[�l�)�>kFI5�n\?W��l��`D ���ʞGbܱ%����:+��a�o?9�Ⱦ�*��t��f��m9�k5����+�xY�l8���V �	g�7g�|U�ƶj�7�u��eHࠣc��9k+d)4y������TH����ͶSTJR�0�}�O��HK�0�ї���k1W��}����|"�f��5�%/F��UxH���N.���w&;W57�#jMu`�w�}XH��Ƀ@�;���Ϊ
g���̛�f�j;�qNuU�W�D���J�R�,�8�Ra����T_]�J��'w }�FS`ِ�����3�m1
#|&�]�$|/�vU��#t�<A�u��\ctd4{�k�nc,1p��f�KM�<�O���H�4�6;�5c����)�fJ^U��4u�)B�LU ːy	����n��q�c|/���#*Z6�뛨��I�E�>�K.2e�ŤJ�ڧt�]��ucV�em�O+��Q�DV�����1�!����Q�iv��q�x9�&k�hOQ.9����j�G{�6�� �~��u�k�W���?~�<d�ާA@9�w�Z�6��Lg ����=N�@-��0��#Ȼ9��%��x��*q�g+Ѥ�:%�*�F��J�Rb�g)�B��J,S�Q��J,Qb��X�ęJ�W�A�3����\%�(1[�z%ꔨU�F�YJT+Q��L%f(1]�iJLU�R�
%�J���%<J�+1Y�IJ�)1Q�	J�Wb��)Q��X%J���h%��(R�P�%���[�<%F*q�#�8E��JS"W��JQb����� %�+�O�%�*�G��Jd+�K��J�P"K�L%2�讄K�t%Ҕp*�P���J�(aW"Y��J$)�E�D%��W"N�X%b��)�D�V%"��P"\�0%,J�*��Y	���B	
Ѯ�A%(��(�_�*��P�'%~T�%���ߔ�^���V�o�ا�^%�V�+%��ėJ�E�/��\�ϔ�T�?+�+�*�R�}%�S�]%�Q�m%�R�M%�P�u%^S�U%^Q�e%^R�E%^P�y%�S�Y%�Q�i%�R�I%�(��+���xT�G�xX���xP��إD�;��_�JlWb�~%Z��)q��*q�[�hQ�n%���]Jܩ�Jܮ�mJܪ�-Jܬ�%nR�F%nP�z%�S�Z%�Q�j%�R�J%�P�r%.S�J\��%J\��EJlV�B%.P�Y��ؤ�F%6(�^	u���#ԱG�c�P���=B{�:�u���#ԱG�c�P���=B{�:�u���#+��?B��:�u���#��G��P���?B��:�u���#��G��P���?B��:�u���#��G��P���?B��:�u���#��G��P���=B{�:�u��#�iG�ӎP��N;B�v�:�u�ۤh���w�����-t���wj��:���n��5�Zʹ�i%�Y��Q����r�eL����SK��s�?5��iә\d>S���"�<��Ls�f3��S
Au��e�a��T�T�4�iכΩiLS�*�*��L�3Ma�0�3Mf��T�4�i�x�qL�1�2���K@%Lc�����L�~{)��o?T�T���y����)��d:�i�<�i8WƔ�4�i�`6�i G�ԟ��a����0�f�f��ԓ�S��d���ݙ\L�:����LݘR�R��L����LI��	�.L��L`�ggS,S�٘���de���p�0γ0�2���N��]�@&&���$ڙE�N����~��'�~f��OL?���A?��&��Ω�1}���}˩o��1�弯��b�_��d��\�sN}ƩO9�g�O�>漏�>d�Lbz��=.�.��az���t�[�.S@o2���י^cz��.�2�K�|���癞�"�2=�Χ��bz�i�\�qN=ƴ��Q�{��av>�� �L��ڸ�NN�ϴ�i;�6b��O�
je�1��t/�=L[�Z���'b��(w1��yw0��tӭL�0�̴��&v#G���zλ��Z�k���
Wq�J�+�.��8��.�K�.f��i3Ӆ\�N53�ϴ�i#�B5h�?a�<�s�	��s���'x@M�l�b�?ah-�����bZ�O����W0-gZ��ȴ�i	�^��1-�'Ԁp�3��|��3��1��zs�fs��zS-��a��T�T�4�iwz:�l�T�t%���y�N��N�y8J9�d�ILe�x7h�?^�a�?^N����sA���}@�q�R���x�D	��0�fg�?~-���T�_*��7����ŠQLn�<���X��ũ�Ꮹ ��4�#��0�\�h�P�4�S	�y���cz�p���ٱ~��6s��r�>|��L��SOփ)�)�)�#G�;��c�s�4��(�n\/�)��Δ���o�J��f���m3A�L	L�LqL�\!�+����de��\2��aL�P�.i�&v�L�`"w{�,����ǁ�Zǯп ����3|� ~~~����ߐ�=���� ���|�����+�%����َϣ�8>>�|���������}�=�]������o�ߴ68ްf:^^�~՚�xxx	�/���u��y�砟�~�:��u��)�Ǔ�َ=���=<��w��(��p�"�C��F.q<�Աhv�?�yۑ�>?�
���"�r���qO�j�ֈ5�������?www �G�q���uno�8�q��7 �C_�X�"�5�u5|WWW ��@�K����'8.
���~����;���yz��\��8���9��ɳγƳ�e�'b��Xc_S�f՚�5�qǆ������jY�9˳ܳ�e��m�k��#<�Z=���ƥ�����Q6�~�B�F[��Q�\�Y�YҲ�C�'.nZ�[l:ŷ���-�m�-�w+�W/�ڊyx�,�Y?�3��;�3�e��>��S�R�ɝ�έ��̝��2�3-��3���S������Sr�=��r���2Ϥ�2τ������-���R��;�S�2�3:��S��S�-ř��dƧ�%d���n�����&����zlt�#Y��UL�*t]���zt��I�;�g���./w��˷]Lq�.=�S�-љ�'Ⱦ%�+/68����`���DWfqt��Np$hE�&���$l ݂2�E��XX��3��Pyvi��&��,���&_�dyu�U�B6��S9��*�E��$�������7Sj~�/u�ׯoْ�_Q�k���6t�Ԅ"�3�4.���O���c�����lӢ�Ett{��F㣣Q���G���C����&/�V=�m�G�/+rbyqt�#B��EL���y��>�����6�O�s����X�4��F�B4�d����%K��_�F��Ӹh��R�\�۵�������o��<�ڵ�V;88h�k�5�j`�8X,���R`	�X, ����<`.0��u@-P���*`&0�L��@�N� ��Lʀ��`<08(�%�`4P�@���@08����P`0 ��~@�����^@O��d@w��i�p ݀T ��@W 	�$	@<�1��� +	D �@`B���F��  �Z�8 ~~��~���� ���=��-���||�����9��)�g��c�#�C��O���{���;���[������k���+���K������s���3���S����	�q�1`7�(��0�� � �hv�;���6��>�>�^�`+��������������� \\\\\\\	\\\������\\ 4�����`=ՎjX��_`����/��ֿ��X��_`����/��ֿ��X��_,��{�� ��{�� ��{�� ��{�� ��{�� ��{�� ��{�� ��{�� ��ֿ��X�k_`��}��/��־��X�k��އ�˭��n��ђ%�fҒf� ���^v��L�y����6�e�(�O��\�kh�A$=F���'����e�O��N
�8���������:y.C*��<�i��s�������R�Qת���Ł��x�"�>D�����F��Co<x��;��2���4��SU���wr�bdΠ�Og�3�7�z�f��C*���i)5�2|-�^HɼEF����k��[h�h5�	\����Yi�W ki���t����\:���m�Mt�o���P�t]��|]|\����%������p9]AW�՘���Gx�2��ҍt�̻��%s��h�K����X�`�xDԸ�c�c�=<�S�y��w��Z�]��9���өƲ�8ʒ�$G�� ��9b$.AX���0���yT~˫���N#s����H����tV�͸�Q��hV7���Ǝ�[���tݎgq�����;�.�������{�'�V��6ڎ'y?�6��[y��o���]� =����N�8���a�x�>N?NO -Kq�)z;�s�<�@/ӓH�d\�A�z�^����U�+���gE�������4�f�O�nG�9�hK�������P�(�r+��v����<TR8(��g����?���=�g�s��oɌ]s��v9�Bi���t�o}��!�┒H�Ŏ	���>�����g	Q��6i֝��y���C6�1%m������8�����K9>�;,g�����?�}�R̰�����I�~vw|�ug�v�l��ln�c�d}wXC�[�܀ Iy��/e����R6�d��_!b�b�Gi���!������!���J��ߠ!CG�t��x��ɴ�_��R�p D[�ʛ2��-9:�b�R�b��ȰM��1�oj���-�=�槗6������k�Ħ&&�Ƅx���o�_
L�\���2-��~u�E3���uK��딴�)�q6SD�-&�٣pځ	)2FJB�:0��j�oZk��tʤ?�q�E�ۿ�i���"�����J�C���ʰɫոFWw�!�{G�q�]�?DFD&���­"�I��H�>ף��]�+��:)�c�P^^^�a99ӧ�t3жo@����D����?;���?4t��9N�
�&Q��2C�'����Q�+=3s�P���K�KO35Z�-��Ȉ3-8��<=<Ε��-,�o�v����eZ%>���h�2顑a┃φY�L�({��e�uKt���HPu�w�Hs7�ic>oK�S�1��lb��m���f5��m��Ö�>(GQ�ȡ4���q�M�^4�����aS0���'!r>1����L�ִ�6���!-.�M���7y��M���08�����Y�'[BI|TH�����r'�w�䴖�c��̖x��U%k��x��+_]�;���n1�&K�%j��E�l�:�撩㖔��wڒb��{f��o�����oZ���=*.96>%.,+'�h�c�W=�nTfNfHL7��[�Lc�%]-G̝��&�0^q6V\<F*.���1�{P��%�G490�[�I�hr`D��G�0�h�?���&2[�唷/�c�`��o��5
���!��,K�PÖglr���3�20c:�劑Ce�x����q�.={vw}yCَA��p_��Ӯ���'9�L�d9N���k��8o�1#��LA����yo�W��59+0O���
�*+Ы�@��ڴwXX�3Ή�%�	��ڔ)vg�W2EffHW�x�eY���/�����9�*�q��ٓi�h��K�Q���kY��o	B̜1=0�c��!�զp���er`�z��b6�r0D�-X;�0��X�M�c�$K�=>�c98/̖�l=��c��ɾ�}�^��ʢs��
��W\`������x�a�vXS�[j(z�-.�kH��-���܀o��=1�:�J�,��e�e��Fil3o����6}5*z9�z&}4���LNJ��`D�tvL�͞g�	;�y�5�l��t��T�{j�7�f'���>RR����H��#Ɇ'�GJ��&ɹa�G��3˝U��gEF):0Jс�':��DF)Z��z� 1�����-�mTg�s��H3��F���jɲl˖|�|���[���I�۹�@n!��pi�-P-��t۟�m�m��N���Pz�ewӿ�xH/�ҊB�C	��=��H���B���H��̙9����{��Qt3�`:����Z�ǎ�G-�[�&� � 	��&�Q41qZ�������2lD�6�˚�n�����l阜S`u:.�[t55f�������2梨[(�g�e�Xͷo�����t����A��������:sˆ-S����c���7p�t�SGm="������N�����{�a� �5����%~���>�����ŜA��*5�k�3�z<ī��U��*y��j^:�ms�s�=�A�q�ٸ9�cY+>�eE�f���cv8���'�w���0�b�x��_�q~q<C=���/�%*�����x���/c<���8�z�8���᭄+�WܤV�����[���`�!�Z��#`a�!z�����Y�c����_��? ��jm|-����}2c��Nb��1���jpL58�{p��⩓�n:�20��G;A�u��%|m�#Zk��(���[VY|ܥS��'0�r{V�����Y�۳��g�O@`Z�u��4�'~V�=�q��*�b�-� �  S��i{�hs�E(O-.Qh����=�5��V,K���a���tUǮB_WgO$t������b���yD��ZQ����AT������p�jN��R}-�\�[Sm�t[
�L�@���t{"���p��˶!-4�ȝ!�> ���"�F�OA%�I�Y��a�,QH���c�z-Q��z�_d�]��uaI�����9�/����Tl;��1$t���?^杕�����*�=V�Kj�{�Ĩ�hQ͎>��}��nQ�nAf��jk���I����I��!Ix�	�.����F/�1d#h�K��H�ɰ�I=�hSŔ�H4d�Y/cP/iOE��I�[��fg4���;�A��O�|f��9��<��iJ�K8���a��>HY8O2J���Dk�C�R
�߮��1���&��Hg�x(r 'x>�~1O��	`"P	_F�vZ��,�(%-PJZ$Ō��֏�a�@�U��U1�UäW�^��ާ�H�a��!8v5c�%�Di5:P�3�jBh(k�Kʲ)�2N�1��+G>����r��3�홍^��]���)Y���w?���x���n�����{����/ߺ�w��➧�]��+����@5=ƺ�a_E�)L�]�ծ�����M�]�!����1�z<���<p91&T��N�<�wܺ�/T
�ʕ&�����Vx���NX��BK�U&���{��-hŀ�\��V�6�m����Vn��l~���Bmi �0�̆���W7��U�M*v�8`�&��!B��T+4��oͰ�ͨ�Ͱ��-� -'cY�g,#@��-A5��PP(��bdw�	���x6ko�������ty>]�N��~@�����Sgepb �yBVO��-]FvQ����z6�����#S����H4)f.m	{�G��t\�zCѮ ��;��7����6��5��la�{�#���_�'�|��X0� ��7�gB�,�(W�_6�sy���!޶���۰��dn����@�*��}��$�+�J%rv^|c�h�s��9;U3w��ש��s���ƓYт�Y
'�I�%�s]0��L&�NqA׹�$�a:�B���q��iQ>O���k�£X3���,'����,��9�S���f�Y�����ӥ�����V�>pW^�yU<>aʛ ���Y�b��k��AY �8rRF��`�'eԮ6\�
pv\mz�4�"i(�Z�CRy��\��k�;�[��ʬ!�j�������Ȏ붏�Zw�E||�M�)��9�KtO�4�jp&G�����~͕��L��A��g�`e�ۼ*ռ��>�q���շ��>�$�2|w���hZٖL���*���`��CH�IY����3P�}d2�BB�xj�3�8��7I ��A�}6n:m|���Q��)2Lr!e[дE�E"�(#=RT}`K�X�;Q��2��_)�|+�EQ���~~D��@ƱY%K���C��C6�CX��*�CD§^�B��(�l�)l�)l�)l�)l�)lO&�laF ��e��	]d�4�Z�$J Ԉ����Yx ,q,�,S����ʢ�ޞCs7]����J+�գ7��iuY- j�Wn~�PW��{�P�R����굷���r}�X,�V,��[Ɲ�3��+�xD�W;�j	w̩�6 5K�=p#k���C�T�F$�Y���tF0������&&�����D�u�t����D��"�MSS�@L�l4C�������!�X�\t�Z
��w�,�R_XO�^X�)˱�1T1d����P�Va�ہ�����H����~v9$�
 hnT&�
�S�%��n���5uxM�	��#U#�:�,O�f� o�����\Y��c�o��P*�ŭ��Xl������nUx���48c�@��H�M�B�����p�Bj-^w��%��{HZy�!�����?/$���w�Nh8w�4��A�a����V���v`�:�,�l|���X���	�������H�<#�B�" �se���
rfQ��K%�2S������ḵ�?l�«��5�5�D�=���=�1���t4n�-�������as5$�i	r~(WRctڈQ"cs)�<�������g!b�H�Y�*l�-����,�q*���Dň�6���������w���/p����������Y���V��yNc��6Nsܑt�z�ɉAg8f�p�_%r�_&~}M1z]��[ӻ��uz�t�	��wT�D���Y��#�9�j�?��EtsD+Hw"������1mޮٮVC`�
w$�3gA 5��������|�}y���R��0��(4}@��!M�@������nO�@�����^GH2s,�	�{��6D5�k����V�Y���8���PA��k����X�ۊ4{$�Ab�#lǭV�z�h������3���R�2ۊ�^((ϜgMg�ʼW}�728�T�l�bR����bU�H�֖�t�h$��X&ÿ�N����,�7K8l�+7��M��P:�'kMO۷fӝ��VW�h�ӯ4v�<x�a�'4y�7�`�dg�����V-_�?j���qմ�]�R��x����&��F�h�c�#:�:�v>��xOp7���x�__WO�W��G�p�d"�ހ�>'INxl�e��N����z�}������	K�GU?l~���u6��h�����w踜hujA��p��D����Չ�=+���+�4�!��	8n��3/�~�O?7`r����)����y�C[�JyC^Zpü��@��PfFE"�>KV����\�4ۊ��2���s�aJ�:'k�-N5C��� /���G�=��(��_���~�O��߷��j�w�Ow*��#�lk��V���o����Uck����,Z��1��p�}�T�}z�x�g��B�q�UF���)�B��c��@1=�:�af8�	��·1��������f��0&���0���2&�(8LL�_�����۠g!l�F�=3�9΅�]�s�`������O�e4�dp��:/��%��ߚ3�o����.������}�����9g4���3��!���ޯ`�β�� �w��[�[T�b����z�|>�4�˲��лx���B-[-`<�ۡz�F1�!a!?�9B���xƌܲ��sL��Q�TWV�-HlX/�EX�����R��ܵ���674O~fu����>�7��&!�ꊱح/ܳb���/�~M�EG�#�L����v���<���fŽ�}Х��W��x�S�r�<����~߰��}�o�Џ Ͱ�6�Ç��a�Tf��C��^BP�,�x�x�4Vx�Ұ�q���/X+�������U���[X�7�ŏ���d��
-�m��%�O�_.n�=�A�XX�	�g:�4��-� ��C߃�{��; �R��/��E�ߧ��6h>ID��Z����~o����W��+����{�i	r�f�R�V�#4��kvK�*��E�½}չlS��.�72V-�Z\a��Ү�r:�"�׎]����o�m^��z!ܚ%~Y�y�w�ۨ�e��j��ƶ,�4�rU��`6LGLf���r:�	�i����jz'y6�,(��k�bq�TI�B-��`�YV9�a�^S8x	"v�F�_rE-Hյ�o�{h�&%p	'U��?��8�Ј��%�^�3\ᆂ�5�u*��V����(`��`��Rۊs�W�i
�=&S��#���F�4>Kx�a��E��x[nc���4��e��hF��Z�����	]MM�A��`�T��#=�)�v��R-;iN�Ém0>T9��^�X:;P�cv�f�L3�����p7����Z��0������D$�W��x��#sou�F͞w�< +M�����~8-0�@��[����"?�<Ҋ�?��aw7U7��@��4�U�aT!��CQe�,W��"�P (�{�2����H�ג�$�:o�EL�7*�A"D���I����"����ʁ��m�<���7�H.808�����Q2«�6R�f�X%�.���@`[/�Eu��������`�����Z��qkh7��Q<��n���[a��X"��T`���������u��n�=�=�e�ڽ�!� �ܗ�����+�?���v�����ݻ��-���W>tmk׮�N� ���JE��O��ͷ�	�w5��=����8^T�(� o�xOF���r8,�2�U\���{������P����l�xW�5a��WZW�;�ߏ�~e�p�Kh�O����"h4�k}̓�/6P� _T`i�*�!�~!{s�����Z>�m��?(�䴢�T�g�q�8r�m+=.�c��iE6�j,����W$)����K��m������ء�}'��|g�h
6��i0�wɋ+���\p��k�mτ���O����� O~��;��f}���JW�k�\���U� �u�z@����)���n�֙zS\h�?�iE����������1��R1;��9X��Qx0�[��dp�?���{�"~�2E�R6f&)���GYk�����1c���a[@.:���u��\���"`Z�c�h��>����I�� 2"���U�	ga����<��m�0W3q��l��u:�WBmqGỎ����". |bw*v�"̳��H��}3 ��g��s���V@��	�X'"�u=�(9�A+ِ�=p4�����x�9�.���"�	���>���O�?L/���8q�u��FS�r�&FC@;s5���jr;x����}U�W�,�7�﵌6�>��f������U�с���.��3YM�E�	yl��H�=QQ���ܙ�13�FN�L"����"�w�F+��!ϻ�: ��X��p:n3R&c���t�����w���l�����7�l����FC��p8}�p��
o@_���\������ �!��0�J���,"-�d�~Bll#,��ȴiڵ@ř"��/`Yy��?jY�|����l���� _��PϦtzcw����'2�#7~aǲ����b������`��Zbg�� ˾�=���f���l���٭ ��8�gڦQ1�~�ڐRBU����/SE���(�=�VI<U�M�~_�x� �@k	z<=�x����|��ң���Fn��ղ0�5_��f���a{QES���X[]�������x������a�
�<]5]��܅d�r�=r$`�K2)��YGKϻ\��LXL�jX݂��^���Jo0.q����*}�����0�9��D���$kx�A3C����dEhA�V1���޸�B��&G9=ܫ�^���M\���<� �V
�IAi�X�9�J�꒎T�	^��,�ģ����H�����oZ,��D*�  �	EM�i_~�e��d�!/S(��Q���H�c>_Ħ����~Oq���Wi&xu᷼�\��:�/��J'�1�\�NI�!�P�?a��`a�P/I���OP5���cN'�Vi��RH�����jڧ�����y'������إ�}�m���� �N���p���;5���;��-���1�VX���?� ���?X(q~�V�� ���_d9���8
�1�� �Sr�'0����^X�`�ΏH�1�� �iJ��Y����G���0MDa%��$�,Ֆ c6㋖*��Z�6���� �(֤�S�LP�2/�4��B��������������JB�1Z�1�����PYm��'3䏑�x�o���ו�"9�����8K� 'Lpf�a�kրE�F�18����s�-�ڠ���R�k�#جE�?�5���S8ր74�vV��`�ăA��f�@�K��%���ђΉ�'�YN�7N�Օ�I�'\Y=g���ʰ� j�&cA�F�6k=oʵ|�K2lWJ��F+<'�<��ä��L�U���PP`��m�e$2cr��>C����nX]�q��8`�_�n߼��gy-Ÿ�ƶ6l���o|�{�˷nU��v��i���gz+z�v�vT�6�jt�h͚F����k^q�^����vu=|�s�n�
k�N�����@�:�ҤN�4�V�#�7���g]�8\\�õ�Ћq8�7�%��.�Ŭ��� �2Gs"2��5��`�f�R�{��6k�����yxbV++�j� �CJ�ֶ��"n�zi�Uػ�	1�͆d��S��M�W��FY��jq�i�����V��Wn�{��ֆ���#��>��cm������"-��X�Z�j�����ǖ�L+���M=�O�������G��&�Cu���O��5b?B�Ǎ�b(SY��SXo�����,�k�B��o*�	.�Op��u_V�����pbF �P�h��pj�>���3�Go��˧�JY��x]Va'eq�������ha+�d�"Cь�����I/�0���6�6�����������n��4a��mkZ���N���2q�$�O�C�;*<����7}�}�&gP2��9�TN~w����p<ĊŪ��5�`7agPֶm���/N�5���s�����&�S�9����:7��;�2-�-D].�#Zr-���ɩ�>�Ŭn��&�9C��F ����Ϥ��.jK`�WΜ9+(sj��񼼳���k!��)G�$j}*��_�.�˥+�dTp�cx�x&��z�1�d�J�)/\ �2;"U�S�7�u��l�HDui�n�wp������'������w��aQ�Gd���}|�+\�|��H�N��Z��B���mG��ʟ[i�������4�d�������<�\ �!�C��k���]�C�/��5��2Cu�)D}ްO�q��jr�yG����ޒf���믨�0�A��,z``�+�����u�H�v��D��x� ���O첁�J�S�j ��$|+�9�5+���}��p��kͶ��XkS���~@q��!!�ɡ4�5�?�>]bz'�����μ��������
p�Z�}C�8!�W@��bd����*������@��@��2����t��%�&��m�����J ���N^��ϑ�^����_��ek�.��߬�kI�ᴼd*<Y��
.4�hvb�g�f�=;�I���a��ӹ,�jO��Kd=$S۞���Q7��"F�F�6��>p����RR���X���Z�g{QQ "YTR�K��&Mϝ9k:- <8�#��2M����.�+\�.���5ڥ��R/b^��</�K��@Fr1> G��
4��SXK����R���+i�����f������O��_��C0���k�����I���&]}�Y�����=���XeW��[��f^_��DE�/ <��89��w����m�FFp�a��{�V��$�7��sL��[��a�)0m��.w��j����(��",��@g5�U ?���`i�H��2�8�JC%�����p-ej�4�4iB0,�D��j�N��4���= ����Qe���E ��:nB<�G�'��y<E�du�%x�,�32:�A��YT�/W�`�/J�<�L>�n|6���+'��Ln���Y���G���Otg����3О�:�2g����G���ԝ}=�	��2}�(�-�ݷOų�XwX�a���X�&�nU�)Ӵ���F��51PW�VC�VC�W#��ƹ���7�|ltj�JH������T�?�T?���"NQ��NQ��K��ͫ��A��{H-�-<�H͗� �j-�����Q��K@w�7e�`2F��־)�%����M�f�?t���M��p�1�ۻkuvjE�g8�$ w5�������-m������j'��i��$"�e���2�Y/y�!�������m=�7|i�x����t3��? �h؆}U�l&(0��t�:�U��.U�T���3�UU�]|1k��aU��M}�H��ߟ3�� ���'~:���!Sp�IVh��epd]$/�ǢP��\2G^NQ�	�^Rfȉ���ꍹ*��XN�1_��1	�[����P����0,E�A��Rju��9.��`H�B?5�y�Y��`�i�e��LU�5���1�۰��&����V8��#�۽k��f#��c���@_mK���!�7�n,Oj������ҋ��Ie�.28���5�a{޼Z�n���657.�v�I�V�C���vU|H�D� ��IRO%k��!0��֦����j�'�P��R�T��p.K��g�~�_�r�x��`R���]~��c��%UԳ$	��hi�Po^5qxM�bF��x������ٛ4{13��6���#;�~�=�i���I��Sܙ�sPh�;�� 6G����Ç<��h���]���o��ȭ���e8]��3@7�i���:�r��}*�+�H*3�)U1"��F��Bu�����{���J����j1���2T/��dxA�h^�D(Q�����`�c� ���֏�����Ky�$/�̏���,G���|��@�f���2@J%B
H�S{=}QF�	:`��g~�%�,b� /Ea�����.���N�Z��΁6��d���Sp��G[J��*%<-������͓�"�R����� ���u׸���)����:𙾾�h�o-o���]4�X:U�������3�!["����9��
)�ȧS�!�RhR\ő{=��ṙ��N'�r�|i�b�*:��r`a7u
����B/|Lw� {�˭Z�,��w�Ѐ���7/�S}@� \�=�|�J5�E �f�{��!	���|��[>-��*��n��͏�5/����j�jn���0-�YJ�
�.Q��MlGm8e��h4/�f@*!�5$e�i~Q�w����{��@ӊ,����#���,�w������od��(�+��ol�����̧?=yd
����ю�q�'�l@,��wL�׮8�Uz|�n�u�����ީ�]�}�W�&rC�vg:W���9�z��"y�i���K��{���}y6�oW^^ܼ��^Aӗ�5%�V/R��K����qt�(\����Xw`0����T���c7 |xI������P��h�#� ��,Cu�y`J��(�H��`O�?־<��L���������[ݺ�[��]�Ӓm,K6`�˶�m ��pH6���$3�>�$�lf��8��d�u�0�yH���k��ل��7a�3��f������,��U�W�w�����~�ABM���6��d��H��S���?]�10=|tҁ���KlM���
�x��^����CS5ߓ�	��t�򗜗R����F�@_���[��Ҕ>��b^O̦V�bo�S�.ÅʇǸtإ��(�
�3��4@)����Q8B��8T*G�����ϞJ�Z�ڍ~�B� ��e�e�D��8��t���퐎g�i�U�Ϋ���M�;3h���;o`��#�*;��Z�����F��I�؍y�KɥU��^b�[
��J`���8Zu�&��F�kBcĶ���t�<�{dk̉�yƼ����̆x�����J:�T(�@Se�4,e(�NarD]�K�W����E�j]���GD��x��vQ���8��tC���o�|��f~Wm�R��|�$�Ѳӎl{"{����×��z���X�O�	`~�&�1p�3[ׂ�R0��\+g�o����1|�%vk����r�#��d<������#[��$��eY��U���L�J�'��?"��g�� ��������?xu�j�)d� ���]Y)=�s����+��_;j`��{'�'' ������f�#�B��"�.I�)�^�{��<�ɚ G=��G<n̕phG�5��&�յʬ�&�%��G�W��;:�z�t؁��S��H��(pq,
����pz2^�{�nq�\)/���L�L((r�HJ7��=�:���׀�|#v������#���RQBN����۟S\�������@͕܎���}�=~km���擓��;��e�����p��[�f�1��W�0�[k���͑�զ�"s��hD����Y�&�װ� �� ��j�eO���3)�B����]ك4�?����g��L��wWZ����<F��+Ms�ݵkp����T���U�Aa�g��#4Г�>��/^�!�&��4�'�w�}�[*���j��_��7NvOFxc#,jL�Ţ5�h��v?o,��C��	p���j~��	m��Rc�.^&]��]䵧��|��)�Js��4�q��8\����`��;�h�/'��E�Z��xH�Y;���V-�l�������%����������Be5�c6;BpZ��w�&��Z�������R�X'�EsM GK�x{#Pn���oHL�h.�}@/Ѧ lm�	��m���ڲ�#��i������u��vu@Bzʥ�[ !o��⯭M�;BC�2�3�BѦ�5Ȋ% q���쿥|# 0e�ښ �)Մ����Z�^�����'Iyh�<��<�a����k,"╊�ɾ�r� �4�!�{C!�k�^my�����c�����*��� ���+ㄶ��r�0,`w�Xĳ%��E�F����.4�Sh����8��	h��@<L���qִ&m$�\1�L�[������ZM˕��s:�~��V��M�_A����=<q[� ���&r\eO�Cg�I�`�f}^��^3��)s�	�z�<2qx��c����s���}vN��׹�Ν:A#T��#�BK���+�1"��}��Ç�7ֶU�y��[�ץ���|`�2� �^RQ[����QKU�ꥣ�8�k�Lth�|�&����FѨ|+4CViW��=F�k����^�k��*�)y/���\]l���-�G�W`/���+,� p+(�0&�WH>,@>�k[zy]�[SX�/.<�=�׋���7�/C��ķ��%��ib�!m5e*�N��Ԃ~�LNV:��}&V�b� x}�<�SQ1~-�&rr�%3tН
�g�(�����T�\�ΌfnK]0u;/1�g�i��HI^#��7�S�׭��}�o����+}�׾��61d��8��S�6 ��>d/������^h\��O�պ�u>D�F���m|E��_�����6Bq�+�\#)	D�19��8���%j��f��W�\�l B#����W�������~�l�;�.,||����6�����\�k���<~}����\!�w�{2Q��X��]��l{���9ۖ]���'��n��;좏�|���۷�=�)�e)5ذcpxi[>R����t8&�vG#��ؚQ)�7w����w�����Y(RJG&���z:�Q]	��/��@l ��(�^�n�ք��2�R��=�\_�0��+�����q���B��7�6�1D��k��@�C��33�ԳBf<O.���$cC`D�����#kŽ�m�)[C�W׋�
O
���X�p-.�V?<V�n�?1^�Ĥ�DeS%!e�W�D<�;�1Yu֢�y<���ܰwro�?l�����?so�LP�;��[�����=C��hΥ���o�e��1���d�X,ihAAQ��|k�b�Y=�PgQ���M��f�I��y:3.7:@�Ȝ����1��#��8*�q8vFMWH׬\Ч��mE��1<'�R%r�s�]>��Z~,eH(��w�D�29�J��`��L�P���
�6t-3z}u
F�z�Z&܄u=8W��V@��j_	�	�؞u�UD×k)��F�q �x�9H�\�c�M�f�BKL9��6���@
~7�Cߧ��P��D?��r�o�`�o�U�7(a�7�66��K�\+M���Ã@�O�W�m�uXJ�A�SKg6�w^ /�x���5@�)�7{Cc�][ �vLe��+���!p��Ax�5C�hL��p�P��F�BJ�Jvaն��&1Zx´�N��濺9�8��)(Jƨ�Ħ=cŝ��M����*^iF��6�\��b���w����$5�w�h-F�ޢ7��Ѱ!�q}�'l���)�S��;�<�k4lL;�#�g	��	���!� ����)T+<S��P9=x�W(���6v�B��Ki	��),��)�R��A�P��_����bfm�\D�SX#�>��ĳH%�	��y"ߞKa~1m �\�^�6E����T��JF�
�B�r^�䏙%J�ۚR�uF��3�_���j"HD�Y�Aa�3�>�y�Ѷ�%��?�?�U<�n��w,�w����:�ʹ�2�'�%9���]y��0��E���0�,#��V�����`�pr���'.�a�Uw��䅖�.��"Ǣ:�«�� l�G��ï4/1�w6���[i�ȭJ��Z��u�uk/
5���r$�	(j%fh��ڰkM�@6�,��&�x�����b^~�fҋ��2�& �SF!�l��Y^����tO�m�O�z9�}�-`$o��༑� W���1+7�nN��]���Y�mర����xUy���3}�̤�EZZ���E<\��t��@�|]�'��qV�A����$q� .犬�X�]���1/bX��X��0��k2\z4���@8��*&?[��1��ff'*��V}M�%Կ�wY�Is>�mی37Ϗ%������?��qq݀����Jή�nZ�jXV�Q[�����O�N!��ԙ�#\�����W(!=�r�Ǝ�Fh9�(�ȏv��6}r�
�a1wC��C�%�"Dy��]L�q�0B�Ѩ��*ɨ�L"��5��_]7ޜ�T� ��ہǟ����i1���@�g�$%V�½i"Ys8���=!�
�q{B5�b������´��=���k��k�߹��̀P&�*�������s����x��[��8x��z���]�������{ �����wJ��vJzԢ��EYSKvP-�G��+�$��K"�f�_r�]�Uvf�]���$	μ�&�5�n�M�/��FJ���X]&Ebrj6�y��ډ6I�ccw���u������V�`W�>,Ym�o���#��u򾧎n�{ϐ�v���e~hϝ(~>��gHݧ�e��iRPMSj�����ܓ�$:� v��)��NQp;Et�=�HU�!哱YH�xܓ�NA�e�=Җ�<g��:��>�%�۶%�	�p�1�
j�Ϣh�Hn8�+^�TI�f��B��Y���D� ��h���o��%��(��
ڏ��N��ɨA�fSQ|�\���Z@��N Ց�*55X�U�$!Ne��I5���)t�Zhig��ֲ�H0��W(�J��y�VGG�@h�5���{t��G+�I�z�kT�TJKv���S���=c1�T�Uz��5�n�zФJ��o�M'f&>6������";��}׼����?/�06;Be�b+B��-�2��!��QCR[҈ �Q0^Q����fѫ~øٸ۸d�1�� N�8�:6�uz}^�@��DۥHo��Q��@Y��H�i~�g{}��^�LEx�my?������Lwl����e[=U��/9Vp�J��͖b��csa~ aU�4���Ts�R�/�m�R���M���������L��H�+����꾮�֚�������sp�P�;���C[	�M� s�x��F��#N�%v��K�g�	��a�6`p��1摽�����c��v�ܷs_y⍹�s�����\vn{���}��_/O�o�9��`ԣ³V��?.���d�KMx�ՄK��_B�+��u�?�	�Bs�3s�p]k_���Zy�����P��!L��9�}`ʈ}��M�k���V��zY���]g��9@�Z_ek��&��#�1�p�<Jǩ���L���d6�v�L��c�[��ܚ�D��Db��5��h��/'J�n�w���l\�)*�����C�m[�I ���;��o��!d?�1�mBF��Vd�I(#��J��t�Z���j6>�L�.A��)��tm�C�p��d���ȷ��RN�R��wU�g�Q��?�����<wa�}T
�~3ހڽ[�mQ2*�=݂i}�D	����������FF
{:��;���Q�/���~qQ�����0{��ғn���+���h0�(sQ̞]w8���Ab~�&��x����s5A^�< �.�#A�֞���urח�F+����Q��9S(��<�m��4]�S-d]���ͭj(meҬ���5�0��$�\
�B���QQ�A(��W�]-���@�Gp�ƙ����כ2@+���S#<��v�pE��)��z	�>2�Jo�$�ڝ�	��n>bAN:9I���h��Q�z*��I��빫�������^��@�0u|Y����Ljz�)�6�����Nm%��~p��w�?�OպyT������|q��/��}c��H:��Y���|����$�Q��M��H�p�Z�_n�>Ե(ڄ�5�e'd?Pq&�譏���o|m��/-ء��&��{*����� �W�Toa��b��t뱃$%����k��n`o>C��8u��QȩŻc0����F�	Y������h��Y��y���coV�����Gc����	Dvf~
���j�{��+���Hx~oI�K�t��Tׄ��7/ք���
b����� ^ �>�pJ�(�K_��ٵU������b��Q�V���{oM��O�pSa�֐%��l�/����HPw�ݻ�(�U�r�� �����E�oA�,��%YD���}x��ox�}�}�}���kVam��u�3�8���L��|�O��}}T��Ex4V�U@���r"Bz��ACy��XD��A_d���jB��ʐ�J�`�4�z�;��� �{[Yl��cq�,�F=6T���s-b�4*tv�*��1q}��Z��x�<��l���]�&����b��N-&�X��K��<�o}�'�=9��6���/Е�I!�O��|h��9S�iG5|�d�`�X�^jY�u�T�	�0ZXhB<�@�n <�H��43s�&���1ʧCK�R�͖�;��mRX|0٦j�޶mz覇����<����5��Fmf5Q�"��b�ԉ���]��v���^����DjX�WKs���=���}�6�3�Q#c�8C���A2$��b�H?��O��d�@� �@e��?����
8��+�A~��Zpb ^h�U�d��K
vW_@+�)����܁�R�sD�dt!�Pc���&gE��f�J�����c$ES�K+�w�e�d��h��*Y]F��R�.�ר��Z�Rk�oR�ԫ��Z��rO��w�Z-�+�wH)5�/������e��|�����@�>X���#{�k$KFd�OF}d�KF=d�M�ed�&��r0C�I�o%�X� ���@�Y?�5��W�H� ?6�T�q��Ev�=�~���%ǳ��Hu�si2���+���oJߖ�6�Om�������b��9�L�anY��!��<#U�c�dZ|����4I����E��4EQ��� ���v�+�sq�����p,1��\l���O��ߢu��חth�oQ�S�Ι��b�]��������+��)�	�Ϥ�~L�/S*s�i�@N+,�&��O�T�nr�`Q�4��
`�J���`�`��R��$�fN 	�_��T0BhٲЦfI;Ѕ�]�N�D��Iq�
jJ���9C�"{4���#��M�#Q�-���F
w�5��A������Zo�����5�C[`CG����jd?��Lc�=#�"�����9���,j٥ej��剘(U��i�Y��cso�	��h�z�i�+z�NF�Պ�irF;�j,��"�k���(�-��rJtC��".Ҏ҉v2���S1��tN���� }U��\UO�f�	1�{���9�fB�$&� )4�D�9
���f�͢�:o��N���ߩb���+ٰ�����ߖ�~w�(��c��֢'�e&5��j�3�Ҡ{'K�l�0pN��bAP?��&R������㢨�gӥSQ���I}��b(-3� ]�,&`rN �01���x��^���\�W���%��t�c�vs�d�V?�%���@���A=�9Xj_ ��z����mN�������1�;T�qb��O�gSX.�ל%`��rG�c�<������Y�#[�R٬��h|����������V}k�]�yT 'g��"�f���48?�zT�/�{�b@D�l��	����\\k��J.o�YHO�����V��3�x�:�~pφ��~�'��QS!�.���j5��H�K��M.�J�u&�1�6[�vO�T��Z���b��� h�E�����ND+���Yr;L	��,	�O�O�
.;�w�f�H	��~�L��qL�i)���W�Ӭ�]��+�,�'��/B|0w!����,�g��bq�LaGg�C}���|�p���W�����*/oN���}H����������G��L$�y�Xd�۟��V6������팃� ���Z���j�IO��e��t��#(
�e6�h�8����1?/����BZ���8��@�kp�ea\�ي���S2E�C���dj��aK*�i�44O
u��LN��F��D�]:�Nm<���a��hT�Mz�Ť�l���}�'�2�=�<x�;�F`Ǻ1v����Yr�2�k�p���)n����E��1���Mx?%p�����U��Ė���,��;#g���xm��?�����+����xD�Zo!�f����s3*�IE�d�Q�h0'2�-٬�k4.wR�0[�|�{��w���,��8�2]�����p�O����q?�'�/����r-�-)��+H��|B �Ȳ@�e�����e��Q�~�Ѧ�wko��gm�&�u�i�7%6��B@�Vꃩ|���Gc���� z@�i,�6S2��mHr���t;�Z�����d���c,O��]^h�����g�n����C�L���@Η��hP�X���I�d����Z���#o.���cB��d���7>-D���k��Z��z�{	�g(����l0�;���4���.�0{Z�Ӵ-?^��*�b�QoRS:�+�鳻=�z�^�O�O��m���v*UJ����$����1I\K�
gtf�1"N��90�m"�<�O���k�r�1����J^S�Gd'��gO������?n�*���h����e�vr���C�\����JS�e,# 8���P�!__�9D��P��!��R�_vB �Ξ+.����t�W�UzJ�x R~RG�\Ȏ	A\*�>���o`�\���gU	=�V�.����w�^�j¤_���3�uQ�#��.w�zh��qě���!'�o�t��5�o��.�@�;��e�s��c���A�3gNٳ|��Ӫm��N�)k�/��p�n|ī�9C�6�?��;]r����FO����z��}^/%sŸ��`���m������$���q䠛� q6ncܦ?�Z�fK�����d�)�i�q�T��ߖ��Թ\56up&,f0������g�4e?�10[�iHk_�e�J�[�d<<��X�뀞R̟Q%v	K/G�<��8�:�%�\�lv����󂣄�����{�m���7��Jwlu]�#f;�{��r�������^o"��Ի?!�"�����N�1>��3	-����磞%��̭�~����o4�� =c!Z�,1��ɵx���q�-��}�$a��=\���Q�U�1V\f�0�`.es�����\�КY��f�L?յ�i�4]�����eDC��O��f��x�s�KT�`�3X���>`��J+���W��R��pm�5ĩ�Y��0su����8�Q��p�L���MNTN���{e�pe����`_���4|b��t���ɀ���x�
��g���TR���kJ�V�W�>��5��-�w��A��=!0ٞ�����2�y-j��e���塞Da)q��B]��1�Z?�	lz;���?-������2Z��=�(\F�5���<���n�h\np��.�����PsG(d+,����\�>0�����+�Sv-���3ۛsG����>Q�j��YacӮ�	��Tl9l�/I�Ъ!��c�SB�-u���F��E;j�����%"8BGaw��\�͚U�#�X�H�a�%�|�'�Ә��%�f���~e��T���C���BKoV��1�43��K�����z�'3��3K�`l�����j�ӆȆlrC�_���o�.�eb�*��fӉ��x�����.�"�[�|��"�[�\�W�;Ԑ�V�X+q�9��q-�G��㪵:�r����:���'ZYZ����X�����N�m� 2z�:;�j�:|&^��;a�SY�I��K�v��?���(ߑ�ُb�T׷2Y뀨 <�����GӋ���`�l���<2}h)yʾ����sETh�8�8{�`_�w=!�cqlPl/,�6��(z㬊��64@�K;�����ÎL:�8c��Ã�^�^�g&� �#�a|�=>@�G� ���>���0��@�T_�-V��p�^�͋�]S_���*5�n�56��1J�����Z-�=��N���z#g4�����v}���6�L)��^?��5�E������zΟ����䶒��&����}���<��g"����6�h����̑֎c�-�J�|򸀛GGzйF�qT ����%���ck׃�tw5��ڢ^@�Z����?��i�4���=�Hf89\-&���og̩a�_9��
 �/&��R3v����Yuf-Ú��;`��Kݱ������/F-�cu	�7d�"�sv��)�I��c��!_r�54�C���I���
l�.!H��o~�G(Ʒ��c'��d֜̇����H8m(�[��EH0؇��O�՜7`ؽuZ��h��b��)�N�)����E��8=���dF?e��L~|�F�7_0�4&$�ߡ�b,�G��U!��8�C*:�d[�j�������x���%�o�3�}K��k�1Qw9B&�����98����_�8Xyo�OHSM#�/�����c�׿[��2� ��䣾�;�����}�9� ��C%���K����"IG�i�Q{�oY��x�!���%����h��>峸JZ�����UM?�0*�m��&9�0E?H)Yc~�֠���@�Q���5j���f��L>�P�i�i�����1J܎���y.��d�Ô4�iТTl�`)H��ҳ��`�]�%�a��p[�F3ԶL�a��!�<����ʇ����-��w�Tв/�Js��
XU�A��K�,�EM��0:-6�QA}��n%��ju����)�Ri�d��-dګ�֟hM�jD�j�'� (�������%�qg�]}Nw�L3��s�it���-KcY�����>0Ll�����B�M��l~�.�$xmɶ�� !D	W�=$$!!���r�k����хaa7�[�u�T��������������dXO��E�P&�m-�L����s}zĐ�ei��0���W�d.r�6E����I�lv��g柱8�[�W
��D��S����)� ЃR�A3�q��8#��U����H���<�8��/Sh�+��D���0��z
`�l�FΒ����}�_Y<�%��w�h@oѻ@��`:5�pH�Qt�Ʉ�(������>Q�B����&����P^��˜Zz��mkc�W^f�ض����GĮxI@�h����}�kӌ*����:\�q�P�N��r�*�.H0�d�J����q=h�8�OE��C%G�O����
�SRwsW��z��:Ȭ�N�����K�]�< Ï�߲�Za�V@��O��O���ҧ蚒p�5�M&)o�M�u(^�`�LIQT-��p�����4¹��CR�i�E-SN��|���^dp�埍[�Ո�H<���Ƨg�-��*;)����Ke�8~7G˸����Q��s޽�=޽���������t��h�ɶ�û�(I�A/qۀ�f�
����Pqص�qX�S\E��㉅�8��1�)���}�X�/�r�R�P��p���X,k����Ū"����<�ԝp�NG�&$ˡ�D�. ˁ:�?�/�(a���oq�������r�����2J�,(��tL�s\��߉7Y��������ip�	T������:���E�P�sE~�D��:E%H�$A+ʋ����H����ܳ��9rC���B���<$Ѝ�[:���E}�
YI�,��XuQ��w4��@H�x�W��ИW6~r{+����]��G<B�KSǅ3��	��0�XP�w��u�"M��<����Vn�ӠwPq�Gw���jh�=�I+[c�pb!��)��Y��j���fFH��{��P�#�����3~Q�g�!�|���S�8NV���JS���H�* I�*(�5�g��A�S�-M�M���	j�CO���OMx���&��������+��.��U�F7�h���'�_9㞢�P�g������T���9�����yۜ�[yy��Q0v�ʯ::W7��`k~uw�2`i�S��lh����u�wD�"� �L$Ra�L������I�C��x�V�T�����-3b
@�d�)*Ѡ޸��s��+GDU�~�P�R!*Bx��S��8~˰\�k`�q{9�\�6�T� �B��sy�/!��l����_�#���~���tJ��8��C�=<����<�l������מ����rND�'��pW�i��"$��������1�ī0�T�c�@�u���x�Ɠu�w�DU�J�Qt:�u ���R���T�*#?:��)'ZȺ���y�I,0�I��auo}Ow������B���*��Hܿ�X󓷪E6���l���B����X�7�$t����.O���,��Kq�����u)"��K�0�M��a�����02�ߌk,�� j7���p��uyl]@����_�F�=��d��%�gX
/��>3��g���ʩ-Kd�>�k�m:�A��p��ve4��Dy-89I-�����\	��g�:Z�����JY}��c�6�=1d���G�^���l�	���f/�<�����#fsQ�V�ѿ]����rGz��dZW��c��w�Vi��'K�^�Ii�)�&s@J�]ϼ����/����,�3�D��5P�ס�	j��ytk��n{q��'qIu|D#�&C%��5Mv�q�]d<�ʻYZ��<=��n_��8=A=q!n˶m�XZ�}a�Aﾊ���gvq��d��}t�O^@�>)���g�K@yo�T��H��Z?P�W)�
�'0�9����7_�99w�8�[��,O�y����˗����<2S�Wg���j�>�"�e?sO�c�K���If�k�vlx�֑y`-��'�Xj�@�"�k��C?�S��i���?~B	J�xP8�*$�����z�_�WK�:4wԅإK�����⠫�r&����c_�������?�6�#�%�a�����ѣ�,����<s��
�������zj+��m�.�nl)�Y�.�4N���=fK�M��Ry�rN��o�U���
	������Yi�)'���J���T�gS�gi���>�M��/���aJsʣ�o8��To��8։����B3R$_aSJX�����a[�=GL��q�|���G�j֩A��B@�֜ K̦�ɸ�h����h��>.���oe����zϩ�
��:F�G�x�#4�:
b�f0|n��1�:��[�&#��J��+`�ȑG�b�?t�O�MGx������#;���|
�lA�Q�r�"Nt����-j���˚{v,m�y o�к6\ٷ������G7:��C�(hQ�x�7��.LTr�xe�$r�KM'�����/�s��o��i#�J%��g��ÒO3���\W5�W58X�Ǹ#���Ӕ�3�3�lEfAZ�.7�Lr˶��(p���r��?ӡZ��Y[���%�<��<�*�K�&��~É"���󬯱==�+������ HD��(����}lhw����-9�z�¾K���k-�Ʃ�,�P�+��,���t]��I��Y��k�Gz�>9T���ٻwM��U�]�m�b��5<�Od�ɞ�ͭ{�@�|��ʧz7�f���R������ފ�?���E���nw�\��0�����f�j*gσ��(͏T�,U7Js��5�9�E���Vi;���æ��_�1���괕Q�9O���ŧRS��-S���E�#�l�G��o�Nx��QYw�8`7�wΛ�����(F�R�T�~�8Y�>f�s8������pXe�X�;�ܧSLŹ�a��
�����zX�-���C�=�9��"oy̽�Qv�#�{�d�q��!|y|��jN�@��^r	[���PD䞅&���q�LG��`Bsz��&ҿ#���LM�)�ʹ�D-�k��{;��ZƖ�Oէ��;�Јl�� ���-j�T�6
̄�X�s�,BV�e��<og6�d�uR�4��='���}��H��K�Ջ.�wɲ&'��d���ttSm����:�`.��^4�(�b(^�phaO0a�S��ež���� ��݀w�6��^Zp�\�YYȬ\�)0��(}�G�֥�?�����ǹ%[����%�~���N�8��G�>��9x����o�T<�v�-k�����O֬9��Z����nq?����΋�7Ix�/�	�ε����Z�o��损���F7��t(��%{�5�n���daS[v�5��PB��ם�t:4B~��x�">)1���c�4v�m�@��+C9@�#@G�y����q'�'�VN@����/���O���9� �<��FgXo�.�h�)w�F髨ԍ��Q�74]�r�Iv�;��:��ɳ�%��E���'��?��]���x���	'��^�o0�x�=�Ey/zI���|�_�>'�����t3�	&�*���~D�]��ל�њ4��m��_�6Q�Ծ���h�[�X��S��ۅ�E�q~�E,:ޛX�b�zӊ@��6��8?�h{Za@!.��'�>�I������^݂\���o?}�����e��Wg��n���k���.��}р��L����dW�J�y�.��R�_��n����xW������Me<h
F�0x��]��ܞ�	

��0���]��v��s@�e��,�}Q۶%�
��,W�m�׹�;�߳�J�0X�h���IOu_}�ƅu8 ��]��U�h����}iT=p��:����x ������;��n.ذ0o˚�d�s<�Ou)Ѱ7��➦u�$������<�e�T-�`󇆄2�&G*9��G��.(Fe��-�.��Rb�t)YV��;0���
��VqFV��������Q �6Gu�˂7f`��R-��Kt+��D�����0���W���e�+��yy���1���wӫd�d9�|TP��īn��VX��.(��tT!{�QT8�ڙ��l�.ls��*b��SH��yx��S�i��1�!�ߓC�r��O<��8�̽��s�`�8��s�A݌����v�PA	�z@��("%��Я�0,�7�	�@����	������"���FOF�<#b��<���Q����s�-�惵sڹ����=���c�#�ze�yt�Gkc86���4J��E�Qu"�`�R)<�)a�1'}��JqbO�^6��5��훭N�ZA�k�S����e�qe��\ �d��bD:Ev��d���Ĉd8�@ e�K�ym�7O���e��Â���5꫎�kgB�\�w�z~��5� �����@�0%1l/��g7�i��m����%�3G�ֹ~o϶۷��7d���$p����5�Q�߅�-w~�⚚��d%�������jE:ز嚅=�}���/����9R����B��LP&L���� ���s�?�-&�G��`&(\�ߢu�`��+6th�q�����Ee3�P�	�2#/Z�첵��eþ��o�6#�e�>�����]ި�*8ǊT�dac�"��ޞ��늞H���\<oϪ�ȵ�y�e9/A�]���*��;�a� h{ԯ�ֽ'@[LP.���χ3|��Ӗd���^����%��d.�j�����`[r3����^)����{b�F���-s�	���eekP"��d&7���t��(B� Jv��,	�c���^�Wlo@TO�f�8Y{v5k{Vgm��풘rGM��)�OY�~�
q~~ީ�[*�/�?�_A��Ex�Ұ��N�Ϊ�H(�R���8>��e�y�Ǫ�j�=M��UX��"����ƈ�)���!̼�y�2�U�,� ��w����m|�>iW��DQ6�}{X�~,�2pF�L�q��I�M��"��S�%B{��8�X���X+�XE|v���v���Ά=z�e0?�%�N�i�avm��˂�[������UI��)����S&��k�8v%�[ly�މ�-��vƂB�e#^�h$�n��n�[
䕦�(`�d�`��)�v��xp��~2d ��%�"������n{$�qs{���]8qW��rv!2,��Q�p�Pđ��b?_S�'G�H��U;�*]Hf>�������1 J��\��0s� ]��]m�H�M���
���6f�MmUx���L(��=�Srk�����2x9�`��Yz���B'v��C��(]��TF�J��0Q�e��eT�$͡4�jB�`�nai�aW�H�V��WO���\N�<W�@{�)��Pq�/���UI�����O�a�G��e��_����5v���&�&��G��?]5�<�'>�V��7����{{г�'ZM4F�;5_�,5wE"S�C9�Ry5jz�e��xk
���)����H�O���_���~	R���л��!E�S��c�&��S*���+�"�)����
H�픍����xp
a��*zIy�7zp��Q����^Ǳȷ���)����q���i�ʡ��FS��n]����#�y.vT9�@h	O��$nbi�W̠��&[���r��Zj�Ћ�t�.Q��(�W�D��U���ǘk(��F�i�W���"|��+B�|&#G֔gΡ�焪A�v�Kղ&s��%��4/)�*����Lr�׫��z/쉹r�\�V:�;"Q�ih����/4�,����^��+~���;޾�.�pݥ�;�����,�	j��<oR��-�-I/jO/Z�ng܁Q��B�r/�.���cOG_���(����C�w���N�[��t�g�$�4Z}�HE�(m0����G��q�w���LҎ�͝����)ie�Q���Лj.8��~y[3`��Ǜd��6&y��p���y����᜵]����"+WT-̇}���NMdůaݫu�E��*�]�u�}]�V��cF\�Kt���p~q���f"�r�s}��c5�ʼ�Fl5��G���1�����M5�hqF�9P���H�f���u�C%��/}�Z�9�Gh�t \p^-�K��Ϟ��w�w#��B����+�Ӽ i�ȗ���K����l/C��?.�s�U��d��
���䛩ޱ�e�8����\b������ۻ:��Y$�>ŧ�t�%���|9\~M8���go��C�h�c{�����#����PY�����BJ�/��&����d��a%(Y����d7�	�b��bz>�֊;��u�-z�%Ɉ��6LP�]4�4=���Q�%��N�MG�@�h�׼}�g�ơ���ѽ����8y�D�	��^ƽc� ߹��ܑY��`�\�|�k�S�w�C�p��y,��|�]>�P8;W�x�翯ѫA���E4B N�y�E�/ �-c��0��a�c�����X���X�17  ���?{�*�߱"db�Ǌ�g
�*>�]R���7\��ъ���5�l�����]�2?վ�=�e��]�"nWK8 ��Q|�"^���j�M�`��U��3�ԟM�.XQ7HЯn�MZ�������~�����@gz` ��`ߒ┳�%�6���Ĳ({_LQ������y�n�"�Fg�zf?�-oɛ3�oY�p1���X~�}�/���>�1�b���Ya�l�MsB@C�j`WO�7_���WwW����=�}�d9��_�4��g#`#�b8)ݺ Ӿ�-�I5G��e�o�-�GD���!]��j ���A���xd��.U�z��qˊ�!y4W�f^E�)q��*��;y��G�NPq�4*�RF���Q��P�~�KG��q�y��/�����3����2��Y(�O�y���q�Sf�2 -�\�����h0�Ϫ�M��Y몡���,7��A?ZXz��F��� ��A�?)��'� ��N��?F�$�o�x�#�<�)&N���ɗ��\�+#�g��^���b�8	��A6ǁ�B���"7���w�'9�7�5B2�`n�ܾ��r2�(
@.<NNt�<#��2�R��!v3��(��S1`��T�K-�.�6PR��}�G���r���^Z\[l��u��U]q��`|�����r�r�����yo�x��������;^W����W^���k/:�t��ֽ��m�m����z���s��Շ�n[ߓ���߶���Bf���U?^?��'�8�������yw���\�
h���-"���dK�����������9�s��^0f�W�y��c�o��>�?�jnlnL�R[��zscc3�Nq}�Tމ�MMiԘ�7���/K[��[8����&<4�K?inn|n����z��k�}���eb �>�А��v�� ����4ߐ����0=N?��l�a�r�~�>���j�#�RfǱQ]4^��J#j5fc�(}�pv�a��Y�Q�+��Gi�5~��qY���X�?�Ȏ���,��fh d���%�)�:�F���S -ս��+o�ܜ�z����U�-�A9���~�3q��H[}�S����Y�8�_k��^��bG2�Nz�QUP��-��ѥ
���x����k�w������(��g@V�_R!�K�sa�+�W��ܘ˥�c�(}��F|�0Ϗ�D&N7V�<&;V,�2�V�v��p�#��5�O֠�KZ��I��R'���h0�vhw_$����$K/�=7�X��2�5�2�(�Cv��qҾ��I�9U���p�m��G�+x��r;<�r�(���Ǆ��������=N�7��!r���"�O�ܿQ-��oP�h��tc��E�(�(�Ҭ4�;�w�,�T~�Yz���x`Xٳǋ�'9������1f!�}*����M��m� �r?�^���ҝ�Kvvuo�u���A��l�t�3͡�@W��o�5ԒK˒�p�eoO]k���)�^�Y�wl���jh4AP�+���Z�eYk~�5�P<�dx�ݜi�3� |׺dǂ�V�}ז��􃤭�Gd��ǽ����:�ГNx7�ṔrJ���g~e��Ѫd��q!��Gu�y��;�q���̓�1��"2'�ox��t���5�����In�8M.s�~���^�2?I��2�e��⯜"�v4��S��>�j���#���}c���d3g�%N�枎��9_��f��L%�A������D0��	Ir>��S�a�T���9����RN��#`��Y(T�p< Ȧ�CK��(��DT<ϔ��:N&���>G��N~#��$��Af�,i*R��q��xzNs��e@��[�6PH�}*��ğ�9�U��]�p	+*�'��ҥ�QTP��3]x���gW]����`��0�*k*IUP���4=��8�:�>�����eE�Ǌs2��5�Z�21�;A���!9j�a�g�J��Z�4c2�D�`pQM����!��*�l���x/;��\�˂��4+�w�~��q���gy�xЧ��Ѧa10��e��W��#�<�+1�
 "��cE���$��;_!���
o�w����ܡ�{d��?��ؿy��]Qv���v6yL�[��e��[�.���yr�DsMB�Z+|ǃ�Xs�b�C����3(���rV��I&�P��S*D�@9�2��Ӆ��.�=�3ӓQ�}-�O��6Pzⁱ�P�*Pt�9��+��,�'�������\]��&(~U1�	��t�������	s �Xm���pX1G��	�J��8�K&륱�ޱ���ig,_�����g�+�9i�!{�4V������#��L{��8u�ĀhI͌���Lہ�q� G�c��sK!Y1sk�;�5Ib��!�Wܼ+��5/�峗�t����u�T�<�V֝�?�^��k��=�L*^���*=����8:�ܹy�/�V�@������T���X&��<��\���	bj�i��]�m+9�e�� ߠ�!�˙�^��^p��GB*̊���5���v����)B�9^y�(vɊ��WW��~;e�Y\��4R���R�*=����V�1� {����$JX���!ձ��A�]�D��M�c���Gp*h�P��hX]���p��s����x҅`�Xc���� !#�v�#W6J?��
ض!��~2q z�f���c���p'�˚�<^���j�H[�Z�p��e&Z����cCU���&�L)d��r��ȟ�֔'~jF�%���f��0E�`�zO�-��0|U�-��TӇ#+D=����?�<'辀�T�8E�5��y&����,���cS�/}�
m���.=��Ss�}^k��Y�^���Q��ļ*��h�ڡa�\ �{o`�s}����m�+�L�z�-S���i�{��7g��݉���.��LSyFM{Kn�ߦ[�j�ސ�+��4P6JЧ�~{{	Z�D�����WU�6�G�/�>��	�F�k^C_+�&>���`��:I�u�m���[�ccS1��:�G`Xml��Q����ua�n�C'�ş>p��a��{���i���{U�����/^�9���_��ǻw-��[��m�n�{џ��Sa*k�W��#H�" ����x`Ǉ��s�us�l��� ����k�u��kn�3����/\�p�(s���5�_�������+�{߫}�b_�6d!(�va��@B���������rU!��l���X��t�,�/��ǉ�x_ӱ�Qp:VOV��=!3g�/�i'+iY����^-9r:�o�u��]�=�?˽�G5E)]�:��}y]E�����ވ����\]��;�-�+4^���l-tQ�?�z�$>����md6��W�l�b�naI���$���X6�5����*�zVa��}^��y��h���}6�HFiu�6$ߔ�f���g�����Y2�yU�G����
��_4�aqC"��#K�8,�t��lG�"�a�������,%��E���̬i�-�Z�qI��B{�Y?S��VV����Vɔ~"��bz�Ĺ$���q�~\�-SSź��+�9��L��:˾��[�Ze��Y��?3kw#8n���J<Y�e�>[�p�58���2듆����$�Y���}��>��)���b�5K��kh��:i���gd���}N�Y�����YԻ#�1����,D�Ϯ"�x����ly|�b۴�����~Q<�xR��?(OJ!_���yG�����(���nP�j��[V賊srKp#���P�e;����Z:�T�v����5�k�?�S��pq�D��n��W�H�=�I��<�0����K�1�]Q�&��>�E�'��HK]���l�)��+˱J�Ҹd�.-(X��+:�YVTT�����%C�da�A�O�W�g��w���kf{
b1�K�$�,�gwIg6�������={\��ץz��b����ᙸ�߁-�/8:�zi�Ώ��	{�"��U�e�'��]ߪ�s�&�����/��R�K"�[ii��z�Œ�a������eSqQy��V;����I}ö��y�[qڴ��9�.���]��8�-~�!W�<#����B^��8;z&�����յi^�]��KEY9��kY��sג�k������;*��-έ;��az�"�/\���lI����ݱeѦ]yEy�����2+6��Z�q�p�IH���Km�0i#����Wq!�*��ӕ�ϬX\QS�`���B_��������c�m�&��Ğy�/_�}U��,�4���PFj[�sd���-�lSE]��C�7��X�֮��J�/�^��d5Cە�[W����j۲����R������sr��ܒ�9�9];:r�s�Wl�(^]��_��]\�o1��f�W4�[j�t�u��~����zt>�X
Y�xq�Ua���ri��j�7>��T���沇���U�Ѹ� Nʥ�������KS�L���M˯[������%J���X�v��勗f�g�o_�S�\�O��$�셟.z�V����ǒ|��m��e�W�/�1�l��Odۍ�����M�ټ��ܼl�������lðNg2�����N�5�@!�d��RAy�X�\:��Y�IaU��e�����gdZ�NVm�ȸ~kY]e�)�`5V8����ZW�X�s�z}�ϯs�d�\���6�������Y�fCv�m�ӵ��նS�K���/&���1W1�t/?�/.��l��y.�f�<ѓ\������g��mu���5�6]���_�K�'"J�˚��Vl�)�^�i,Y�yY���M�L���e���JY�a:MPo���|`p������]�K��Y8�,s�8���Ґ���hܔ��đ������c2�dY�unߟ!���/�ɓ����r9���P�i�-��~D�����3s�=�Nڐ�[P�(�ҏ�F������7�e�����&��t2���,�~(Ê��C�_:���\>�{��z�&}U��6i���d޺�5y���:�ˡ����kO~�(�X�Tez�A��u���I35X�ţ~a�9*~G]�qȿ���ﯔ����+)-�]����#21�#b�Z.�+o����!��l�� �:I�$�]�\� }LwP#}��w��d�W%�����LU�m�,Â�tA��V�O�s��_�2�3&�hVP���!ǖ8}��O�ѯem���b��Dw��h�*t.�\ng�nK�oʯZ�>TP���q:&�h�U�����%O�N�N��-�]�f��ٽ��sK���ȕ�<x%�p�pUX����*�J����I��|Z#�ZN�]Ao8ߨ}a�{�<�����>����^אB�����߽�a�˂6>��M?�9"h��-;���?t�K�o>m}z���ȵ�aE�f�o�ӗ��q{�M�5=м���-w��~Ǯ���j�k}��Pۓ;��|bW������'���#�ю�gS���.Mi�3�	F]�U�u�nX
:z�W���m��q�yAz��8N���8���ͫSoɟ����<��&���W��G��S������������{Sh�K���{��r�����f
}��վ���~��&��/����|�Ty��^h��חBa��xOx?�D�N�_7-���t�������9Ë8-^5\7�e��k��ÿ�W_�o���MeiJS�Ҕ�4���[T��a�e��NgFZF^y)P
�@�28����4�)MiJS�Ҕ��jNS�Ҕ�4�)MiJӟ�>���Gn��wA�w�_����
NMiJS�Ҕ�4�)MiJS�Ҕ�4��]О4��.�����*�G沢��-2��^ce�d�Q�2Y�{^-���I���eCR����A-��u�[ղ�(�q�l�N��[�^�gղ�\g�����&gى1�;��)�R-Sb,p�e�cjY&��T˺�1zb+��Z6$�ɖԲ���רe3q���-�+>�JV�N-�H^Q�Z���j9�,��P���R�>��΢,pe��(���Eِ�.pe��(�EY�,�gQ8��=�P٤��_ 
YC���lDi7�	� ��{�D�ֈR����->��=�RH7چ�0�"���O/F�� F�I+J�h��	n^��%�xI!��||G��~���$
��ss�5���NR��U�m U|}78�0V��n��xx�au�NԆ��zG!_$�O/�}\�U��8(d;���a�n�B���OP�Tᫌ������=��a�2�Q5�üm7i�L��n��|���`M�� UT���
o�p�� �f���?
)|�
�\���Í��
}�|E��W7�1^�P;�R��!��Q�s�����C*R�k��$�p�<\� _%���ƭ2�揣���Um��:	,"�+"��V��Y,��k������R��e��*xF8R		؊!���[!��{�a�s�T#���Q^p[k~-0�;T���~>2!q�F�1>Oh}�j���\���p�8�j�&�y_@�d���K�{��^nk湡�6B�!uL���ܣ�BX�H�Jn�#,FR��2�����u�j�]���Xϕ�j�Z�U=G��������kpOd��� �W��!կC���s�����o-��W�q�!��T�([��+d�� �,
b�j3�pl�̑+��Z����q�^�ls�n�.0ָ
�~.�`�K+�൐�F�����m�����4�8��h���h-/x��͢��c�ƅT�H��!�k@���W��՜����5��s94+ϷXT�!�'|E�`\��k�bW��F��GħX�*��|D=�q��xZ����>i~S"�Ğ�;K%ƯL�����Tl��C�?G��<)��|��|��$� �D�"NZ��O|��<⾪����)^%�AP}Z��(����>�Ss���F�y�����,P-��E�/�T1��Ořeu;ϗ^U턡����U�2n^ ��j~��	������D���gVu��!4�Z_���}�r�J5z�"qФy7��5�J�<��4��7�M�I�q:�H»�i�Ӽ���\W<r"Igao�^u-���ݫ��au����\4��Y�c�W!��#V�s���y��$v����/`�8Bn�;�ͧ��5V=�Y;�eM�3}�4ᾩ�xuۢܓ����+�0H�CH��k�Gw5�腳[ռ�a?������ɕ8�%�&�i6�"������$	��/?���VH��e�;�hܖɹDذF�x�G�?.�ש�t�&��B��&էH�8���v�v�Q~w)��&I0�_ٚ	\n�O��}�|,2� �@��6�dqq;����|��v���3m�X(��Ί�\!lկ��뾊E�q�#�K����+�|�T���V��{;Ij��[v�6�)Ȣ��ًZZ�в#z���R��>Ԋq{�'xt��<ǵ��Ym�w���L��5�������w��?��qlF#Z����;x�u`���hS�D!i/ڕ���R��5�v����jox�q~L~�~/w��lQ%m�1Όg#$j�5ֺ?�0�����u�vpZ�/ti����U]�8��^��و��Jh��1h��$�k��.H���@o/�!:1��k���kV1cڶ�ZB+a�F�C�aЄ�n|�c��_�,�I�R������~�k#G��ׄ5y��ۊ�V����z�_u��f>��k����Bz�;��I����m�eѼZy�\��=���ą���1ar��W�g���5�ڍ�n�'��Jc0
��Q_0P�4��J�oh8Q��o��w�����{�*�!o��Xȫ���G��?8��(�`�X��Pgg�����P�t���a���=�Ѻ38PZG"l��a_D�'����~����+�ĢJ$8�x&�Qwث��a%:�Uv��*�>�7�nQ"^����x�hU�O�b��5�Q���nt�}�a[í���p	��A���L9�+����߫��X��P��`f`  ��p�Zi�*�^wt4�(a/��E��'R�DF�����̦�����XFG�a��x��AD	��������Qe�*����U|%ʰ�d�X+8����8c�P�;�d�ao����"�����(L*�f� r�]¾C��QFClpBK��~�����[�F�Z�y<��0󆫻�C�~w8�W���73X�1��^S�}4����Ç�ܤq��!��	B����n�T�#+aEeG8�G���暚��'R=�ͬƄ��Pp(��q����P��zܑ�` �cTb��h(���qX_�r 8
Ď)�p�(sV�̀���Qo�2����� �����f�G|�(���Zi���7��Vd+T]�;�``��b�xs��m����3�$�Q,�x������� <�ҷR�E�ppx'iE��a�H4�����~������a�K%a9���=���[@ς:0+�FC�^�&3���RE^���� >'þ~_��'{/D�ha"�PW)��d�B3B���@�Q�a_�;�sW�C5�V���Ss�J�����f�$�P���:������� tb� ��Hl��4ɠLI�v{3N��^̂c��*e0���B�8���
�t%؏d`��y����ڵ`�#����f��8C�
D�"���@��qL�V�Q3��Vr�x6vXpϳ�9�ݪTwc�k�~�T��x��N�x1�X.���^Hh
E�y��u�(�kT��@񈗥�`�'2�UE�%EШHs!�G�AG�� ��rA�P.�M^OTs����|<�6G;�M�p�(��}jOQ�"�l?���D�;I�0[>�3�`����N �xkmVz:[z�5t7+m=JWw�޶��&eEC�+��}m���{z��n��=�t�(�]mMUJ�������[i����֌�����=Mm;���щ}�����
[Pe���Ø�n�nlE�a{[{[�*������l�������qO{C�ҵ������7�mG[GK7Vi���ы-�mJ�^T��ֆ�v�T�H���k��:�ݶ��Wi�lojF��fHְ��Y,���vW)M�v4�Y���͇���km�MX�_��m�L��Ύ�nT��ewo|꾶��*��������	�N���L0��YpaP+)�V��Ӝ������z�������c��c�w�m���_���u>�K?H?H?H?���ӏRh������ �)�k@��Br'Y�Կ�'�߅�/�����*m6�1��Z���l���Z�gf��е�w8�x�ĵ���b���u|N������÷��f�BRLJ�Ȗ��<�U�05�=d+�jRi3Gº���$_ ��SH���})���T��{���ڨD�h&]J���zZF�h%�]�M� �����	��A� ���#��-�%z�~��EBO�_�I���$�'�:%�3�R:#��/I.zN�-��˻%��G
�������;d�t���N�U�_�MzD����k�%�u����O�9�u�-���2А�i~*.r���C�������(py�������g��Mr��K.p).U�e3pi.=��p��c���壨}�<
\^ .�.? .������tR�p).����4�N��^�2\F����]��^�rp�py��\�\�'p�9p��<'S�-9��
�P����%	�������	\n.���1��A��i��%��p�p�!p���&��]� �j�R\v����\n.1�r
��p�"py��\������#���"�ѓR9�Kr�S�6���.^�r3p��L����C��i�2\~ \�p�%p�W9,��Y�M^$\^-�Z^/�.7�o�������p.�Rq17	�"�R	\6 ����Cl���{���˳�����e#.�a�\J��z��	\��r��..�.��3���2\^.�iPʤ��b��l.;���2\��%\>\>\��<\�\�\f�˜�G&�>�_Γ�r	p�.k���r�x�K��\&��g��C��i�2����cI�,.�������.� ���ˣ��z~N�Q����� tp�\n.c��o��W�����e��*p�p�����K*�7J��Oj�~� p9\��{�˧��C����e�r�����Nɔ��3茼��$;�9�%�w�� p.�/�) ���y��,p�p�!py��N���t��]��{]5���T\����K)p�\��a��n��.�������M��f�*�r=p9\������)��=��/��f���b���I��� �Ja�r��\._.�.���ғ�D�s�)y)����O�.���\�Q�r
�|
�<\�\~\~\~#��Qٯ3�a]�|�n�|�n��q]��k�~�u�O~C�~�rpy�<\���9�o���r8*+�������dM�pM�Lj2�M��51gҡg.�W,���66�b��h��+�p��2Qj��ԋ�ѫ�9���,�ӟ���O�9g�>��G?z������gnbb�-�*F^�����M�\�c�Ϥ'&�E\��Sn|������JL��	e�k���S =�hmu:[[OpF]]��AO�9������'��5�CL�o7�!�Ǉ&.�bc&1霮9�0�`��싅 ����7���X��&Y!�S\�Xl����ӓ)@L�`y�O��K
^�긘T����f0
M&�L�Y�ZB�)�c֨#F���ٰџ6�A/�0���<���A>� �>�tM��\.��~��l�̄�0�p��\�%K��b�� ���(Fq�1����&�á0^��qp��H`Ī�r�x����2������t}�9xx%4V�+^	�LT�ή���N"&�5�r�d�bϊ��D\��<<S=�/fj�����}�Q�<5:��d��4�\������G4���i�j�a�S�1������79�:tČ�X(@4fW�]"B�:jF��!b��G�?#,���#<�]���Đ�A�,5�q��&��0�J`��	׵8�b�GI
*�@5PP�E/�^&�֝UK ����&�bj7�۸��Fj6�o��l�g5��s�O\�V����]��ټ�����ؤK�%��l�A�\0[��6��~�������l�f˙�����;�� ��o��]`n��
b�xm�ͅb[!��l$f�%�zŅ�q��g�;C�!a"f+5�Y@}H��) e6ݾ}��¥K������p���,0ϲ���Ϝ�Dg�a]bg��.�N=��SQ��ٖy1;n��>Y.�4�3��a�X
O���T�+f�/�� �詅�����	���1��m��s<I	₨�5�N�e���ϰ8fUUv�?�uԨ\��Y��s8fY��k�89?�
3�X4!��b�6��\��e�,"����5aI�`���,l�,T�h�pmY(8�I��H�j����t'�l7������:��]����
oaq�K���$.�_j*To�,]���=�������u�ɄX��D,�U?��sj��1k1<,���'y�4Q�yk���a+�Z.��8�}�"w��Z^�X��ϵ�w�~�:�ͻ�g�����]�X��>�7Շ�s��DÇ��K�3�X���jW�\4�"H-F�!��q�j�cT#���a�K*�se��2ㄢ�~�`��O+�V�>���u��V���J�W���O�p�Z����5��V51�<�����!k�S+_�Y+��$������:���_:h�T�jA�`�
�H��m�L�Ia�7%�V\+\�^���x�r����&z1^Jj�-��Q&6�:�n����2�{V�Zl�5eTr�n�A8W�e5Q���-$u��X�r�N��w^����X��D��Ĭfj�.&}1x�n�'�[LxW�Q.'9�|'b\�U�Ԛ9U8Ux��t�d�d+;�a��4n�\�b�A����	�8�v!K	�|a�U�j���� b>^1?��;ѝ&��H�IQKr6��2(�+��2�m ��8�nv�d��v�.��0"i��'&��gh��z��� ����,���>�r'�{%\�[Xo�f���������L��0~|��q���h��˖��L��fJ�'l�ڒ-3Y�)�٩�D�m��;k��'	^״�b�>D�1�x�255��� T�ȹ� n:Lޖhɂ��idk�pD�`bq�`��-~Dd�pB���D%v+F�SF��،��%5g����2����%���KZ��Y�fdY����kRu�K�>v �X�Hԑ8$	>�Bݖ������e�pebOdj7�3�(��a��5�d�E�jc����۰����f�6�b����$�C�bb�P���ƽ�T�u&6�D��]b����R��ǧ/��\��K��������L𼜼��M�}R�۔T�dˠ6�l�l�\�+U�����h?w�쩗NMۦm������+S�A�@3�����L٬�f_LnVШo��)hlg���g�V��d�Ls�!�,jgb\�����ٱ���ܘ�Dl�˅�k�����F�a�ڌ�a����l�Ԗu�p�0}������s�ϯ�_?V�,tr1������m��6�;��Fe [��}����֙�o�����Dx��iv����%�r��~ז!�?���A͙ص��n�k����]�S/�m��[1���KLO�%j�MM���l�;��8׬�H�f�;s�����s�fԉI��F͙����9�B�.�������z[R�k�2����~Е���jK�[���̬�Sc�0aH����V�8�6��v�C�����b��)���'�>R?W�W��o�ݘ�l�-9	⢭��	��h�${RD G���)��`�쀣^��NŰ��n�g�	jYF�a�hx2���)��z�X�j���9y#/������s��N�q���y����U v��Po@��qMp�|������嘁0�i'Cz�����a�eKN�ie�1K���V�[���ruD���rC��_�4�GUJ㱰�J���a���(�w0T)��h�ݍ�2P.�K?���B�ҏ;�K��`����;߲S�tz�����Qku��U�T�'N���� ��7HTw��y��*���e�Rϩ���M����۬����I�t���oy��O����/ܻ����a��[N��q�릝��C�e�JRND�����ž0x�i�K��8�r1�=:C����6Ǚ�*��>wd���gk4���#��@m����Xr�|�`m�s1�s
����Ꞩ{$�t568�
�띛�j7�۸�� �������HfwZY�5G�����v�s���}!�v���f���cs˺5W�mذa�Ɔ�k�9��JԨG�)�9N+��z"��L�v�4N)��uɢ�9Q����L�h8Q9�������Z���/�<e���߳�4�߇?]�ȡ���O}b��~�h��+��á�ްc2H"��xg����gߗdoc�.ˇ�dI֩(���$���K�ȒߌJ������w}\��y�9s�������������C�]��<�3V�T�cr��Ԋ9��q8���M*��E&bxZ���6�U|�L�<E��mA�TΥ���h���?�8IAR�av�M�l�v�P�����	�K�c�=�������Z|�&=&��$dh�l���p�?/!�"V$�(��~����x���hRV���4�M M�-���w�d��.�'�.7٦�>�Sx��x����|$��"x fI� 4��Ə��8���I�$�[�`r�}1�Bh� *V���:
���g�}�Ѽ��hr@�F�:�
(�(�ȇ�~���r������	{U�[���m����&bP	�|0�'�8&&w��*��w ���6���߯������(v��R��{���?9$.%��8oV󕢧���ؚ<�Ύ��G��2�D;�����}{�y�F�[ �	?iL�У�v�0yOn�>M'M�Ӌ����W�� t��P�JCsr��V4�O*y���u̚� N��5� t�'�#�����o^б�r	�y��D�%�9ȭw���+UV��k������"��ĥ��W-�R�%�]Es�Rf	!��ΉP�s��G^Cl�	�O�f�1E8zt�΁�lPo�*��?���
]��=r�qIgi@�046����#7�����i���`h�ʿB\ �W�g<�nkǤ��_D��Xl�4|��D Q8`~������W����O����"�j�Z	�҃�w8��xE�m��GE�(T�w[F
���L�ߺT̈�즫��RXlO��aX�F��➻� ��I;����$m�4��:f�.<*��!�T*O(77�i�ݾ�?]H��{]��Ax�i��-�w�[ƽqT���$,���*=!Q������Z_6P��Bo[x���ķ'��λt_%����V��ө��O <c|d�ҍη&S�>��3^/�=�<Е� ��U*�&
����-ly8U�]!�ܦ����A�KP���l�Y�K_�K7ʬF:�T�Ct�=`���C�Y_gmIu+4��6�`��" ������E �k#
Y�Y��Y�!E�EO!�mE���V������(P��vF���1�{n��|��N��d(��,���c �ů%�? ���S��!
�0��!
������_��b'�� `L,�{w�E�A8�4�Æ-Z���y����7w�Կlz�����n��"�˶�ɝ4�dˣ�\Mx����:����E�>k����[��;���(����tz9����㡢�^���8#�V�r�.�'�H�b�2��8����1N�i{�HI؞!�z�{Hb�.Z@����:�������@ 9O�|"D2E�Pُ5�K%EG�!�v;�	�T�9����.�wme���z�5����)^O-pkr�|���ع�TLR��)IzҤs�SH�WnL_���k�A�"�"A՜JU�ֳ�l.�g����t�?��s_����T���َl���A���j6�7~�V�gpN����{��J˛�.���Uֺą��{�^(���۱}�&I8s)���.���g)7��)���Wwδ�I>	H��x�Ӓ�����!�n�b���!�j8+��3��Cq�	��\��p[rV�5���YO��E�C��*�g��k?$u�ӯ9�4���~a�"uڈv,bšM�H�{��E\C]�/Rr�m�?���yu�7#X�*�V4�B��O�sk�O��D�����ق���b�?��E��b`���7�~𦎇�<1�u�w���c���v��r���; �p��  �!w|���C��g�V�+%�\r�����jO�f�*}:B��F���Z�7�tt��^2�r�	�ĲT3�c�e�b�R$�'2H�Zdc� [x��{z�������ͬ�]�[�ψz-�{+d y�]sx��FA�"�w�K�y'LS_�t�o�9>p�02����s̨+�}��j]7�����J8*��G9��o��_���}-:�HE��]���Jg�"��C(,W��*Զ��e�������d�����k��p�r�SF�)����g��&���^�Y�"���q� \̿C|���K��a >�7M�a�� ��_�98��"��<wր5��� �M6���ks��_�'�"��&W%��T��{(���*
� F�rds�ä�y\|Ќ=MK����wH� @� ��?11�{�~���Ø��@E���ʝ��[�7�4@[T	�>o�F
-y�p1��O��f]c��`�j����4�-7J��` �ݩ�_��]�L6��u�*M��R�h�$N��:�j~���/pw>����s��δ��'�I�:Z���.�^�5�b7�۵��ͤhR���&	��{�*�p	^/��O��k�бb��k�j�-jD_m��o\��L"s�_׋y���33#�"��J�p恽�_`��m��L�$�;bj�o�Zs��ep���Y?�8�ƈ\#��}&����t����[��5��Y)9|I��Ĝ7Q���C�+�:�e�������9J��,�^�y����J=|��� 5%6K����Ѵ̮������GW|�3�͜z�+�%"s}���Bo+�Qz�F!\���iwư>���d��K���L3�ܫ貹믇�/Ӻ�TQ�_��I�{��a@�"t�1�ao�Y�bX<��8}Ey���#��r�S�[��"�S8�Y��٠����-�,)�>��ch�.�$�x�ߥ�,�o_
pN�#�*F �W���'�##�cdC�}�S�&���yƂ�Q;�X� c��s%k[^���A��H
u�������eN�̛hݮ���(?��JzrD��� ɚhK~E��K\�E� ��+I��\˳�o�;Z�e�V󵖿.�-$*�b�u�o��w��A)0[B��-Wm>���)q��v�8m�K�^�Ḩ�w[a��r�gۜ%8��,�@�{�HCԯ!Ibu{�ׄ�Q݀+/�k��t�����lB��U�N����1����[�0���/4j����x�ƕ��*O�җ��A� �Y��U��������YC��?���d�֫��^����nI�u���K�=UL�ԳK��e��E��KV��\ʙ����/�U%u��J��=4x�:�iN�����ę��FZ7Q��O��Ί�ϳ*����]��nn�
��ekTHk_m�7�]RW�J��-�f��T�O6��/.,��*sA�
�.;������}exìя��ݲ[+W_�Y��kr�mDj����ɟ�7��������%5C�*"��fi�O��S�qM���9��e�v��B�~��/��7P�!�'�qt��eq�������i0<^����BQ�9k�`�Uܰ�P5s�sTÔ���>��x-�Y�K@��ؗ9�C2�h�dN���_��gc'�	F�I@p��"�p��@��p`��ߥY��0�����+������8{�:�`b�Q�����״ܯ��Z���.|�<�;���11�*sX+H�����v`� I9:a��&�r�/�4����'�����-�K��q�x�bq��ӰM#�p��.4�r���� i�>:U��32�:��.S�0'
��1�%�M��>���d݀^.���}��V�i����Y�G����K���q1R�a$rr7IM�y����;�#�[/���^6Sι�;�AV�ƅJU'� Y'�`lE�N���?5ͺ�,F����Qi�L��a�my#Q�yN����97G�N39�VG:�{U{����/�pI"����$Mh�qW�=�/��Μ��o5ױke�9�
��\��M�xR��]1���2%�.����҇������ڛG' c�d\+�vK���f)�8�
���"U%�� �^��ʌ)y�����Y���K�Y�>dm6�T��&}��D�hU�Ь�>o˷v�I����w�e����17�����A�,��G́��ĕR۷zn�7�Fd�7�P�o�y��kJ����\����X��H��8R !w� ��_ׯ�x9�܆%�o &�~���Nn�X��c�m7I������`�1�z�����t���[H��^O�/�����I��Al��z'�1���$GW�za��,N�a���@-Z�@
N�X槨g�("D.B�BמMH'�z.5���˔�=�`'S �v
OTt}�h�:�s\�����U��[�}�ÿ�ۭ�~�9����34[�i��'���a�=����%�̋���~Կ�a�P�ɤ�I���BʖB״3�M�v�g���Q��"�\T���'^v��Ĳ�/����b%�(q�疺BĈE�)��x0)�x���9�ȹ��'%�]�dΠ�:ǛG�8�U�L��r�`.Lx��c���H05���}h^���_�i;�Is��0$I~�1a?h����?8>F��?&@��|�x�W�"G�{�#C����R&,V�Ы�HC\zc��"q�
� w������ʥ���9��"����Xvg���� �4��SvTů�ʯи-H����X%ʕ�ZW9�G�$�q��WN�c�_�LB`��p�0�
�j�cgʅ�h�Q�i�ٿb5*�X�;:4���2cc���T�S[���w|���<���fI6OwF�����y�F�|�hl]I�"4S�ˍs���7_�熆I/C�e���k_q��.�i
!О8�Qb�V�Z-o�^�)��������0��]
endstream
endobj
223 0 obj
<</Type/Metadata/Subtype/XML/Length 3056>>
stream
<?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?><x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="3.1-701">
<rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
<rdf:Description rdf:about=""  xmlns:pdf="http://ns.adobe.com/pdf/1.3/">
<pdf:Producer>Microsoft® Word 2016</pdf:Producer></rdf:Description>
<rdf:Description rdf:about=""  xmlns:dc="http://purl.org/dc/elements/1.1/">
<dc:creator><rdf:Seq><rdf:li>BiServ</rdf:li></rdf:Seq></dc:creator></rdf:Description>
<rdf:Description rdf:about=""  xmlns:xmp="http://ns.adobe.com/xap/1.0/">
<xmp:CreatorTool>Microsoft® Word 2016</xmp:CreatorTool><xmp:CreateDate>2026-01-07T15:20:52+01:00</xmp:CreateDate><xmp:ModifyDate>2026-01-07T15:20:52+01:00</xmp:ModifyDate></rdf:Description>
<rdf:Description rdf:about=""  xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/">
<xmpMM:DocumentID>uuid:DF5BECBB-AC68-4935-AA47-42401E6639C6</xmpMM:DocumentID><xmpMM:InstanceID>uuid:DF5BECBB-AC68-4935-AA47-42401E6639C6</xmpMM:InstanceID></rdf:Description>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
</rdf:RDF></x:xmpmeta><?xpacket end="w"?>
endstream
endobj
224 0 obj
<</DisplayDocTitle true>>
endobj
225 0 obj
<</Type/XRef/Size 225/W[ 1 4 2] /Root 1 0 R/Info 13 0 R/ID[<BBEC5BDF68AC3549AA4742401E6639C6><BBEC5BDF68AC3549AA4742401E6639C6>] /Filter/FlateDecode/Length 441>>
stream
x�5��VVЃH�`aww`c؊݁؍�����-vv������{����5k������;*���/��+$�gH�ܐ�l�Jl~H\NH|^H͔ (y�|�g|�W|D1�;�9����BIG	ĠJ�ʢ�#�Xġ2*���
P�P�Q�PuPQ���M��$$���Z�Z�5ڡ-:�=:�3:���+z�;z�/z�7�` ��?c !C0#0�1#1
c1���q�ɘ�I��)������HC:f`fa6�`.20����K��+�
��k���؊,l�fl�>l�v��N��n��^E6�� �rpGp�p����8�<����9��<.�".�2
pWq�q7� �Q�;��{���x�Gx�'x�gx�x�Wx�7(����H�&��A��>$S�g%�%*5#$�0� 
t
endstream
endobj
xref
0 226
0000000014 65535 f
0000000017 00000 n
0000000165 00000 n
0000000228 00000 n
0000000501 00000 n
0000003304 00000 n
0000003478 00000 n
0000003723 00000 n
0000003776 00000 n
0000003829 00000 n
0000003999 00000 n
0000004240 00000 n
0000004506 00000 n
0000006987 00000 n
0000000015 65535 f
0000000016 65535 f
0000000017 65535 f
0000000018 65535 f
0000000019 65535 f
0000000020 65535 f
0000000021 65535 f
0000000022 65535 f
0000000023 65535 f
0000000024 65535 f
0000000025 65535 f
0000000026 65535 f
0000000027 65535 f
0000000028 65535 f
0000000029 65535 f
0000000030 65535 f
0000000031 65535 f
0000000032 65535 f
0000000033 65535 f
0000000034 65535 f
0000000035 65535 f
0000000036 65535 f
0000000037 65535 f
0000000038 65535 f
0000000039 65535 f
0000000040 65535 f
0000000041 65535 f
0000000042 65535 f
0000000043 65535 f
0000000044 65535 f
0000000045 65535 f
0000000046 65535 f
0000000047 65535 f
0000000048 65535 f
0000000049 65535 f
0000000050 65535 f
0000000051 65535 f
0000000052 65535 f
0000000053 65535 f
0000000054 65535 f
0000000055 65535 f
0000000056 65535 f
0000000057 65535 f
0000000058 65535 f
0000000059 65535 f
0000000060 65535 f
0000000061 65535 f
0000000062 65535 f
0000000063 65535 f
0000000064 65535 f
0000000065 65535 f
0000000066 65535 f
0000000067 65535 f
0000000068 65535 f
0000000069 65535 f
0000000070 65535 f
0000000071 65535 f
0000000072 65535 f
0000000073 65535 f
0000000074 65535 f
0000000075 65535 f
0000000076 65535 f
0000000077 65535 f
0000000078 65535 f
0000000079 65535 f
0000000080 65535 f
0000000081 65535 f
0000000082 65535 f
0000000083 65535 f
0000000084 65535 f
0000000085 65535 f
0000000086 65535 f
0000000087 65535 f
0000000088 65535 f
0000000089 65535 f
0000000090 65535 f
0000000091 65535 f
0000000092 65535 f
0000000093 65535 f
0000000094 65535 f
0000000095 65535 f
0000000096 65535 f
0000000097 65535 f
0000000098 65535 f
0000000099 65535 f
0000000100 65535 f
0000000101 65535 f
0000000102 65535 f
0000000103 65535 f
0000000104 65535 f
0000000105 65535 f
0000000106 65535 f
0000000107 65535 f
0000000108 65535 f
0000000109 65535 f
0000000110 65535 f
0000000111 65535 f
0000000112 65535 f
0000000113 65535 f
0000000114 65535 f
0000000115 65535 f
0000000116 65535 f
0000000117 65535 f
0000000118 65535 f
0000000119 65535 f
0000000120 65535 f
0000000121 65535 f
0000000122 65535 f
0000000123 65535 f
0000000124 65535 f
0000000125 65535 f
0000000126 65535 f
0000000127 65535 f
0000000128 65535 f
0000000129 65535 f
0000000130 65535 f
0000000131 65535 f
0000000132 65535 f
0000000133 65535 f
0000000134 65535 f
0000000135 65535 f
0000000136 65535 f
0000000137 65535 f
0000000138 65535 f
0000000139 65535 f
0000000140 65535 f
0000000141 65535 f
0000000142 65535 f
0000000143 65535 f
0000000144 65535 f
0000000145 65535 f
0000000146 65535 f
0000000147 65535 f
0000000148 65535 f
0000000149 65535 f
0000000150 65535 f
0000000151 65535 f
0000000152 65535 f
0000000153 65535 f
0000000154 65535 f
0000000155 65535 f
0000000156 65535 f
0000000157 65535 f
0000000158 65535 f
0000000159 65535 f
0000000160 65535 f
0000000161 65535 f
0000000162 65535 f
0000000163 65535 f
0000000164 65535 f
0000000165 65535 f
0000000166 65535 f
0000000167 65535 f
0000000168 65535 f
0000000169 65535 f
0000000170 65535 f
0000000171 65535 f
0000000172 65535 f
0000000173 65535 f
0000000174 65535 f
0000000175 65535 f
0000000176 65535 f
0000000177 65535 f
0000000178 65535 f
0000000179 65535 f
0000000180 65535 f
0000000181 65535 f
0000000182 65535 f
0000000183 65535 f
0000000184 65535 f
0000000185 65535 f
0000000186 65535 f
0000000187 65535 f
0000000188 65535 f
0000000189 65535 f
0000000190 65535 f
0000000191 65535 f
0000000192 65535 f
0000000193 65535 f
0000000194 65535 f
0000000195 65535 f
0000000196 65535 f
0000000197 65535 f
0000000198 65535 f
0000000199 65535 f
0000000200 65535 f
0000000201 65535 f
0000000202 65535 f
0000000203 65535 f
0000000204 65535 f
0000000205 65535 f
0000000206 65535 f
0000000207 65535 f
0000000208 65535 f
0000000209 65535 f
0000000210 65535 f
0000000211 65535 f
0000000212 65535 f
0000000213 65535 f
0000000214 65535 f
0000000215 65535 f
0000000216 65535 f
0000000217 65535 f
0000000218 65535 f
0000000000 65535 f
0000010080 00000 n
0000010292 00000 n
0000031720 00000 n
0000032046 00000 n
0000086890 00000 n
0000090030 00000 n
0000090076 00000 n
trailer
<</Size 226/Root 1 0 R/Info 13 0 R/ID[<BBEC5BDF68AC3549AA4742401E6639C6><BBEC5BDF68AC3549AA4742401E6639C6>] >>
startxref
90720
%%EOF
xref
0 0
trailer
<</Size 226/Root 1 0 R/Info 13 0 R/ID[<BBEC5BDF68AC3549AA4742401E6639C6><BBEC5BDF68AC3549AA4742401E6639C6>] /Prev 90720/XRefStm 90076>>
startxref
95399
%%EOF